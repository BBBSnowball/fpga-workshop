
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

package pcmdata is
  type tSAMPLES is array(integer range <>) of signed(7 downto 0);
  constant pcmsamples : tSAMPLES(0 to 46817) := (

    to_signed(-30, 8),
    to_signed(-30, 8),
    to_signed(-32, 8),
    to_signed(-37, 8),
    to_signed(-42, 8),
    to_signed(-43, 8),
    to_signed(-37, 8),
    to_signed(-28, 8),
    to_signed(-18, 8),
    to_signed(-9, 8),
    to_signed(-6, 8),
    to_signed(-7, 8),
    to_signed(-11, 8),
    to_signed(-14, 8),
    to_signed(-18, 8),
    to_signed(-24, 8),
    to_signed(-31, 8),
    to_signed(-36, 8),
    to_signed(-36, 8),
    to_signed(-34, 8),
    to_signed(-33, 8),
    to_signed(-31, 8),
    to_signed(-28, 8),
    to_signed(-25, 8),
    to_signed(-27, 8),
    to_signed(-34, 8),
    to_signed(-41, 8),
    to_signed(-44, 8),
    to_signed(-44, 8),
    to_signed(-42, 8),
    to_signed(-40, 8),
    to_signed(-37, 8),
    to_signed(-33, 8),
    to_signed(-29, 8),
    to_signed(-27, 8),
    to_signed(-25, 8),
    to_signed(-22, 8),
    to_signed(-22, 8),
    to_signed(-26, 8),
    to_signed(-33, 8),
    to_signed(-37, 8),
    to_signed(-36, 8),
    to_signed(-31, 8),
    to_signed(-24, 8),
    to_signed(-16, 8),
    to_signed(-8, 8),
    to_signed(0, 8),
    to_signed(5, 8),
    to_signed(7, 8),
    to_signed(5, 8),
    to_signed(-1, 8),
    to_signed(-10, 8),
    to_signed(-17, 8),
    to_signed(-19, 8),
    to_signed(-16, 8),
    to_signed(-12, 8),
    to_signed(-8, 8),
    to_signed(-6, 8),
    to_signed(-4, 8),
    to_signed(-3, 8),
    to_signed(-3, 8),
    to_signed(-3, 8),
    to_signed(-4, 8),
    to_signed(-6, 8),
    to_signed(-10, 8),
    to_signed(-10, 8),
    to_signed(-5, 8),
    to_signed(4, 8),
    to_signed(11, 8),
    to_signed(14, 8),
    to_signed(12, 8),
    to_signed(8, 8),
    to_signed(4, 8),
    to_signed(0, 8),
    to_signed(-3, 8),
    to_signed(-5, 8),
    to_signed(-3, 8),
    to_signed(2, 8),
    to_signed(8, 8),
    to_signed(12, 8),
    to_signed(16, 8),
    to_signed(20, 8),
    to_signed(21, 8),
    to_signed(21, 8),
    to_signed(21, 8),
    to_signed(23, 8),
    to_signed(25, 8),
    to_signed(24, 8),
    to_signed(23, 8),
    to_signed(24, 8),
    to_signed(24, 8),
    to_signed(21, 8),
    to_signed(18, 8),
    to_signed(18, 8),
    to_signed(17, 8),
    to_signed(14, 8),
    to_signed(11, 8),
    to_signed(10, 8),
    to_signed(12, 8),
    to_signed(13, 8),
    to_signed(13, 8),
    to_signed(11, 8),
    to_signed(11, 8),
    to_signed(12, 8),
    to_signed(14, 8),
    to_signed(13, 8),
    to_signed(12, 8),
    to_signed(12, 8),
    to_signed(13, 8),
    to_signed(12, 8),
    to_signed(11, 8),
    to_signed(11, 8),
    to_signed(14, 8),
    to_signed(16, 8),
    to_signed(15, 8),
    to_signed(9, 8),
    to_signed(5, 8),
    to_signed(5, 8),
    to_signed(7, 8),
    to_signed(11, 8),
    to_signed(16, 8),
    to_signed(22, 8),
    to_signed(27, 8),
    to_signed(29, 8),
    to_signed(30, 8),
    to_signed(29, 8),
    to_signed(27, 8),
    to_signed(22, 8),
    to_signed(16, 8),
    to_signed(11, 8),
    to_signed(10, 8),
    to_signed(11, 8),
    to_signed(13, 8),
    to_signed(16, 8),
    to_signed(16, 8),
    to_signed(15, 8),
    to_signed(12, 8),
    to_signed(8, 8),
    to_signed(3, 8),
    to_signed(2, 8),
    to_signed(3, 8),
    to_signed(3, 8),
    to_signed(2, 8),
    to_signed(2, 8),
    to_signed(5, 8),
    to_signed(8, 8),
    to_signed(6, 8),
    to_signed(1, 8),
    to_signed(-3, 8),
    to_signed(-6, 8),
    to_signed(-6, 8),
    to_signed(-5, 8),
    to_signed(-3, 8),
    to_signed(-1, 8),
    to_signed(-1, 8),
    to_signed(0, 8),
    to_signed(-1, 8),
    to_signed(-3, 8),
    to_signed(-5, 8),
    to_signed(-6, 8),
    to_signed(-4, 8),
    to_signed(-1, 8),
    to_signed(1, 8),
    to_signed(3, 8),
    to_signed(4, 8),
    to_signed(3, 8),
    to_signed(1, 8),
    to_signed(-4, 8),
    to_signed(-13, 8),
    to_signed(-22, 8),
    to_signed(-26, 8),
    to_signed(-22, 8),
    to_signed(-16, 8),
    to_signed(-10, 8),
    to_signed(-8, 8),
    to_signed(-6, 8),
    to_signed(-4, 8),
    to_signed(-3, 8),
    to_signed(-4, 8),
    to_signed(-6, 8),
    to_signed(-11, 8),
    to_signed(-17, 8),
    to_signed(-20, 8),
    to_signed(-17, 8),
    to_signed(-9, 8),
    to_signed(-2, 8),
    to_signed(2, 8),
    to_signed(3, 8),
    to_signed(4, 8),
    to_signed(4, 8),
    to_signed(4, 8),
    to_signed(3, 8),
    to_signed(1, 8),
    to_signed(1, 8),
    to_signed(4, 8),
    to_signed(10, 8),
    to_signed(14, 8),
    to_signed(17, 8),
    to_signed(20, 8),
    to_signed(23, 8),
    to_signed(22, 8),
    to_signed(18, 8),
    to_signed(13, 8),
    to_signed(9, 8),
    to_signed(4, 8),
    to_signed(0, 8),
    to_signed(0, 8),
    to_signed(4, 8),
    to_signed(8, 8),
    to_signed(9, 8),
    to_signed(11, 8),
    to_signed(14, 8),
    to_signed(16, 8),
    to_signed(15, 8),
    to_signed(12, 8),
    to_signed(11, 8),
    to_signed(10, 8),
    to_signed(9, 8),
    to_signed(7, 8),
    to_signed(9, 8),
    to_signed(13, 8),
    to_signed(17, 8),
    to_signed(15, 8),
    to_signed(10, 8),
    to_signed(5, 8),
    to_signed(4, 8),
    to_signed(3, 8),
    to_signed(1, 8),
    to_signed(-1, 8),
    to_signed(0, 8),
    to_signed(6, 8),
    to_signed(9, 8),
    to_signed(9, 8),
    to_signed(11, 8),
    to_signed(16, 8),
    to_signed(23, 8),
    to_signed(24, 8),
    to_signed(22, 8),
    to_signed(20, 8),
    to_signed(21, 8),
    to_signed(19, 8),
    to_signed(13, 8),
    to_signed(5, 8),
    to_signed(1, 8),
    to_signed(1, 8),
    to_signed(3, 8),
    to_signed(3, 8),
    to_signed(3, 8),
    to_signed(3, 8),
    to_signed(3, 8),
    to_signed(4, 8),
    to_signed(5, 8),
    to_signed(6, 8),
    to_signed(5, 8),
    to_signed(0, 8),
    to_signed(-5, 8),
    to_signed(-4, 8),
    to_signed(0, 8),
    to_signed(2, 8),
    to_signed(-1, 8),
    to_signed(-3, 8),
    to_signed(-1, 8),
    to_signed(3, 8),
    to_signed(3, 8),
    to_signed(0, 8),
    to_signed(-1, 8),
    to_signed(0, 8),
    to_signed(0, 8),
    to_signed(0, 8),
    to_signed(2, 8),
    to_signed(6, 8),
    to_signed(9, 8),
    to_signed(11, 8),
    to_signed(12, 8),
    to_signed(13, 8),
    to_signed(11, 8),
    to_signed(7, 8),
    to_signed(3, 8),
    to_signed(0, 8),
    to_signed(-2, 8),
    to_signed(-4, 8),
    to_signed(-6, 8),
    to_signed(-6, 8),
    to_signed(-5, 8),
    to_signed(-5, 8),
    to_signed(-6, 8),
    to_signed(-10, 8),
    to_signed(-14, 8),
    to_signed(-17, 8),
    to_signed(-18, 8),
    to_signed(-18, 8),
    to_signed(-16, 8),
    to_signed(-12, 8),
    to_signed(-10, 8),
    to_signed(-11, 8),
    to_signed(-13, 8),
    to_signed(-15, 8),
    to_signed(-16, 8),
    to_signed(-19, 8),
    to_signed(-23, 8),
    to_signed(-26, 8),
    to_signed(-25, 8),
    to_signed(-21, 8),
    to_signed(-17, 8),
    to_signed(-15, 8),
    to_signed(-14, 8),
    to_signed(-12, 8),
    to_signed(-10, 8),
    to_signed(-9, 8),
    to_signed(-7, 8),
    to_signed(-5, 8),
    to_signed(-4, 8),
    to_signed(-6, 8),
    to_signed(-10, 8),
    to_signed(-11, 8),
    to_signed(-9, 8),
    to_signed(-7, 8),
    to_signed(-8, 8),
    to_signed(-10, 8),
    to_signed(-11, 8),
    to_signed(-10, 8),
    to_signed(-11, 8),
    to_signed(-13, 8),
    to_signed(-15, 8),
    to_signed(-13, 8),
    to_signed(-9, 8),
    to_signed(-5, 8),
    to_signed(-3, 8),
    to_signed(-4, 8),
    to_signed(-6, 8),
    to_signed(-9, 8),
    to_signed(-11, 8),
    to_signed(-15, 8),
    to_signed(-17, 8),
    to_signed(-17, 8),
    to_signed(-15, 8),
    to_signed(-13, 8),
    to_signed(-12, 8),
    to_signed(-10, 8),
    to_signed(-6, 8),
    to_signed(-2, 8),
    to_signed(1, 8),
    to_signed(1, 8),
    to_signed(0, 8),
    to_signed(0, 8),
    to_signed(0, 8),
    to_signed(4, 8),
    to_signed(10, 8),
    to_signed(16, 8),
    to_signed(21, 8),
    to_signed(25, 8),
    to_signed(28, 8),
    to_signed(29, 8),
    to_signed(27, 8),
    to_signed(23, 8),
    to_signed(20, 8),
    to_signed(19, 8),
    to_signed(18, 8),
    to_signed(17, 8),
    to_signed(17, 8),
    to_signed(18, 8),
    to_signed(19, 8),
    to_signed(18, 8),
    to_signed(17, 8),
    to_signed(16, 8),
    to_signed(16, 8),
    to_signed(16, 8),
    to_signed(14, 8),
    to_signed(9, 8),
    to_signed(3, 8),
    to_signed(-5, 8),
    to_signed(-14, 8),
    to_signed(-18, 8),
    to_signed(-15, 8),
    to_signed(-9, 8),
    to_signed(-6, 8),
    to_signed(-6, 8),
    to_signed(-4, 8),
    to_signed(0, 8),
    to_signed(2, 8),
    to_signed(-1, 8),
    to_signed(-5, 8),
    to_signed(-6, 8),
    to_signed(-4, 8),
    to_signed(-2, 8),
    to_signed(2, 8),
    to_signed(8, 8),
    to_signed(16, 8),
    to_signed(22, 8),
    to_signed(23, 8),
    to_signed(20, 8),
    to_signed(16, 8),
    to_signed(14, 8),
    to_signed(12, 8),
    to_signed(9, 8),
    to_signed(3, 8),
    to_signed(-3, 8),
    to_signed(-4, 8),
    to_signed(1, 8),
    to_signed(9, 8),
    to_signed(14, 8),
    to_signed(13, 8),
    to_signed(6, 8),
    to_signed(-3, 8),
    to_signed(-9, 8),
    to_signed(-12, 8),
    to_signed(-16, 8),
    to_signed(-22, 8),
    to_signed(-27, 8),
    to_signed(-28, 8),
    to_signed(-25, 8),
    to_signed(-21, 8),
    to_signed(-18, 8),
    to_signed(-16, 8),
    to_signed(-16, 8),
    to_signed(-18, 8),
    to_signed(-20, 8),
    to_signed(-20, 8),
    to_signed(-15, 8),
    to_signed(-8, 8),
    to_signed(-1, 8),
    to_signed(7, 8),
    to_signed(15, 8),
    to_signed(22, 8),
    to_signed(25, 8),
    to_signed(24, 8),
    to_signed(19, 8),
    to_signed(15, 8),
    to_signed(11, 8),
    to_signed(9, 8),
    to_signed(8, 8),
    to_signed(9, 8),
    to_signed(12, 8),
    to_signed(15, 8),
    to_signed(15, 8),
    to_signed(12, 8),
    to_signed(7, 8),
    to_signed(3, 8),
    to_signed(-1, 8),
    to_signed(-4, 8),
    to_signed(-8, 8),
    to_signed(-13, 8),
    to_signed(-17, 8),
    to_signed(-21, 8),
    to_signed(-23, 8),
    to_signed(-23, 8),
    to_signed(-22, 8),
    to_signed(-20, 8),
    to_signed(-20, 8),
    to_signed(-22, 8),
    to_signed(-24, 8),
    to_signed(-25, 8),
    to_signed(-26, 8),
    to_signed(-27, 8),
    to_signed(-28, 8),
    to_signed(-25, 8),
    to_signed(-19, 8),
    to_signed(-12, 8),
    to_signed(-5, 8),
    to_signed(0, 8),
    to_signed(4, 8),
    to_signed(5, 8),
    to_signed(4, 8),
    to_signed(3, 8),
    to_signed(0, 8),
    to_signed(-3, 8),
    to_signed(-7, 8),
    to_signed(-12, 8),
    to_signed(-13, 8),
    to_signed(-10, 8),
    to_signed(-5, 8),
    to_signed(0, 8),
    to_signed(4, 8),
    to_signed(5, 8),
    to_signed(1, 8),
    to_signed(-8, 8),
    to_signed(-19, 8),
    to_signed(-26, 8),
    to_signed(-28, 8),
    to_signed(-28, 8),
    to_signed(-30, 8),
    to_signed(-33, 8),
    to_signed(-35, 8),
    to_signed(-33, 8),
    to_signed(-27, 8),
    to_signed(-18, 8),
    to_signed(-11, 8),
    to_signed(-7, 8),
    to_signed(-7, 8),
    to_signed(-8, 8),
    to_signed(-9, 8),
    to_signed(-10, 8),
    to_signed(-10, 8),
    to_signed(-6, 8),
    to_signed(4, 8),
    to_signed(17, 8),
    to_signed(28, 8),
    to_signed(35, 8),
    to_signed(38, 8),
    to_signed(39, 8),
    to_signed(36, 8),
    to_signed(29, 8),
    to_signed(21, 8),
    to_signed(16, 8),
    to_signed(13, 8),
    to_signed(13, 8),
    to_signed(15, 8),
    to_signed(17, 8),
    to_signed(19, 8),
    to_signed(21, 8),
    to_signed(22, 8),
    to_signed(18, 8),
    to_signed(9, 8),
    to_signed(-3, 8),
    to_signed(-13, 8),
    to_signed(-19, 8),
    to_signed(-24, 8),
    to_signed(-26, 8),
    to_signed(-24, 8),
    to_signed(-22, 8),
    to_signed(-21, 8),
    to_signed(-21, 8),
    to_signed(-20, 8),
    to_signed(-19, 8),
    to_signed(-17, 8),
    to_signed(-18, 8),
    to_signed(-20, 8),
    to_signed(-24, 8),
    to_signed(-26, 8),
    to_signed(-25, 8),
    to_signed(-19, 8),
    to_signed(-8, 8),
    to_signed(4, 8),
    to_signed(12, 8),
    to_signed(14, 8),
    to_signed(13, 8),
    to_signed(13, 8),
    to_signed(15, 8),
    to_signed(14, 8),
    to_signed(8, 8),
    to_signed(-1, 8),
    to_signed(-8, 8),
    to_signed(-13, 8),
    to_signed(-12, 8),
    to_signed(-8, 8),
    to_signed(0, 8),
    to_signed(8, 8),
    to_signed(12, 8),
    to_signed(8, 8),
    to_signed(0, 8),
    to_signed(-9, 8),
    to_signed(-15, 8),
    to_signed(-18, 8),
    to_signed(-22, 8),
    to_signed(-26, 8),
    to_signed(-28, 8),
    to_signed(-27, 8),
    to_signed(-22, 8),
    to_signed(-15, 8),
    to_signed(-8, 8),
    to_signed(-2, 8),
    to_signed(1, 8),
    to_signed(3, 8),
    to_signed(4, 8),
    to_signed(2, 8),
    to_signed(-3, 8),
    to_signed(-5, 8),
    to_signed(-1, 8),
    to_signed(10, 8),
    to_signed(23, 8),
    to_signed(31, 8),
    to_signed(38, 8),
    to_signed(44, 8),
    to_signed(50, 8),
    to_signed(50, 8),
    to_signed(44, 8),
    to_signed(33, 8),
    to_signed(22, 8),
    to_signed(12, 8),
    to_signed(4, 8),
    to_signed(4, 8),
    to_signed(12, 8),
    to_signed(23, 8),
    to_signed(32, 8),
    to_signed(34, 8),
    to_signed(31, 8),
    to_signed(26, 8),
    to_signed(22, 8),
    to_signed(17, 8),
    to_signed(9, 8),
    to_signed(-3, 8),
    to_signed(-15, 8),
    to_signed(-21, 8),
    to_signed(-18, 8),
    to_signed(-9, 8),
    to_signed(1, 8),
    to_signed(5, 8),
    to_signed(2, 8),
    to_signed(-2, 8),
    to_signed(-3, 8),
    to_signed(-1, 8),
    to_signed(2, 8),
    to_signed(2, 8),
    to_signed(-3, 8),
    to_signed(-11, 8),
    to_signed(-17, 8),
    to_signed(-16, 8),
    to_signed(-8, 8),
    to_signed(2, 8),
    to_signed(10, 8),
    to_signed(15, 8),
    to_signed(15, 8),
    to_signed(12, 8),
    to_signed(9, 8),
    to_signed(9, 8),
    to_signed(9, 8),
    to_signed(3, 8),
    to_signed(-7, 8),
    to_signed(-15, 8),
    to_signed(-16, 8),
    to_signed(-13, 8),
    to_signed(-8, 8),
    to_signed(-5, 8),
    to_signed(-1, 8),
    to_signed(4, 8),
    to_signed(7, 8),
    to_signed(6, 8),
    to_signed(-1, 8),
    to_signed(-12, 8),
    to_signed(-25, 8),
    to_signed(-33, 8),
    to_signed(-34, 8),
    to_signed(-28, 8),
    to_signed(-20, 8),
    to_signed(-14, 8),
    to_signed(-9, 8),
    to_signed(-5, 8),
    to_signed(0, 8),
    to_signed(6, 8),
    to_signed(7, 8),
    to_signed(2, 8),
    to_signed(-5, 8),
    to_signed(-8, 8),
    to_signed(-6, 8),
    to_signed(0, 8),
    to_signed(10, 8),
    to_signed(23, 8),
    to_signed(37, 8),
    to_signed(44, 8),
    to_signed(42, 8),
    to_signed(32, 8),
    to_signed(21, 8),
    to_signed(10, 8),
    to_signed(5, 8),
    to_signed(7, 8),
    to_signed(15, 8),
    to_signed(24, 8),
    to_signed(26, 8),
    to_signed(23, 8),
    to_signed(21, 8),
    to_signed(23, 8),
    to_signed(26, 8),
    to_signed(20, 8),
    to_signed(7, 8),
    to_signed(-7, 8),
    to_signed(-16, 8),
    to_signed(-18, 8),
    to_signed(-17, 8),
    to_signed(-16, 8),
    to_signed(-18, 8),
    to_signed(-22, 8),
    to_signed(-29, 8),
    to_signed(-32, 8),
    to_signed(-29, 8),
    to_signed(-23, 8),
    to_signed(-18, 8),
    to_signed(-15, 8),
    to_signed(-14, 8),
    to_signed(-12, 8),
    to_signed(-10, 8),
    to_signed(-12, 8),
    to_signed(-15, 8),
    to_signed(-16, 8),
    to_signed(-12, 8),
    to_signed(-4, 8),
    to_signed(4, 8),
    to_signed(13, 8),
    to_signed(21, 8),
    to_signed(27, 8),
    to_signed(28, 8),
    to_signed(24, 8),
    to_signed(15, 8),
    to_signed(4, 8),
    to_signed(-4, 8),
    to_signed(-10, 8),
    to_signed(-13, 8),
    to_signed(-11, 8),
    to_signed(-6, 8),
    to_signed(1, 8),
    to_signed(7, 8),
    to_signed(10, 8),
    to_signed(6, 8),
    to_signed(-6, 8),
    to_signed(-23, 8),
    to_signed(-38, 8),
    to_signed(-45, 8),
    to_signed(-44, 8),
    to_signed(-41, 8),
    to_signed(-38, 8),
    to_signed(-33, 8),
    to_signed(-23, 8),
    to_signed(-10, 8),
    to_signed(0, 8),
    to_signed(3, 8),
    to_signed(-1, 8),
    to_signed(-6, 8),
    to_signed(-6, 8),
    to_signed(0, 8),
    to_signed(7, 8),
    to_signed(13, 8),
    to_signed(19, 8),
    to_signed(28, 8),
    to_signed(41, 8),
    to_signed(52, 8),
    to_signed(54, 8),
    to_signed(51, 8),
    to_signed(48, 8),
    to_signed(48, 8),
    to_signed(47, 8),
    to_signed(44, 8),
    to_signed(40, 8),
    to_signed(39, 8),
    to_signed(39, 8),
    to_signed(38, 8),
    to_signed(37, 8),
    to_signed(37, 8),
    to_signed(36, 8),
    to_signed(30, 8),
    to_signed(19, 8),
    to_signed(5, 8),
    to_signed(-8, 8),
    to_signed(-19, 8),
    to_signed(-23, 8),
    to_signed(-22, 8),
    to_signed(-18, 8),
    to_signed(-16, 8),
    to_signed(-20, 8),
    to_signed(-25, 8),
    to_signed(-28, 8),
    to_signed(-27, 8),
    to_signed(-22, 8),
    to_signed(-15, 8),
    to_signed(-10, 8),
    to_signed(-7, 8),
    to_signed(-7, 8),
    to_signed(-8, 8),
    to_signed(-9, 8),
    to_signed(-4, 8),
    to_signed(4, 8),
    to_signed(14, 8),
    to_signed(21, 8),
    to_signed(25, 8),
    to_signed(28, 8),
    to_signed(29, 8),
    to_signed(27, 8),
    to_signed(19, 8),
    to_signed(9, 8),
    to_signed(-1, 8),
    to_signed(-10, 8),
    to_signed(-17, 8),
    to_signed(-21, 8),
    to_signed(-21, 8),
    to_signed(-18, 8),
    to_signed(-16, 8),
    to_signed(-20, 8),
    to_signed(-30, 8),
    to_signed(-42, 8),
    to_signed(-52, 8),
    to_signed(-57, 8),
    to_signed(-61, 8),
    to_signed(-64, 8),
    to_signed(-68, 8),
    to_signed(-71, 8),
    to_signed(-67, 8),
    to_signed(-56, 8),
    to_signed(-39, 8),
    to_signed(-27, 8),
    to_signed(-24, 8),
    to_signed(-26, 8),
    to_signed(-25, 8),
    to_signed(-21, 8),
    to_signed(-16, 8),
    to_signed(-12, 8),
    to_signed(-8, 8),
    to_signed(2, 8),
    to_signed(15, 8),
    to_signed(26, 8),
    to_signed(32, 8),
    to_signed(33, 8),
    to_signed(32, 8),
    to_signed(31, 8),
    to_signed(29, 8),
    to_signed(27, 8),
    to_signed(24, 8),
    to_signed(23, 8),
    to_signed(23, 8),
    to_signed(26, 8),
    to_signed(30, 8),
    to_signed(33, 8),
    to_signed(34, 8),
    to_signed(28, 8),
    to_signed(17, 8),
    to_signed(3, 8),
    to_signed(-11, 8),
    to_signed(-19, 8),
    to_signed(-21, 8),
    to_signed(-19, 8),
    to_signed(-15, 8),
    to_signed(-13, 8),
    to_signed(-13, 8),
    to_signed(-14, 8),
    to_signed(-16, 8),
    to_signed(-19, 8),
    to_signed(-20, 8),
    to_signed(-19, 8),
    to_signed(-17, 8),
    to_signed(-15, 8),
    to_signed(-14, 8),
    to_signed(-12, 8),
    to_signed(-6, 8),
    to_signed(0, 8),
    to_signed(6, 8),
    to_signed(12, 8),
    to_signed(17, 8),
    to_signed(22, 8),
    to_signed(27, 8),
    to_signed(30, 8),
    to_signed(29, 8),
    to_signed(25, 8),
    to_signed(17, 8),
    to_signed(9, 8),
    to_signed(3, 8),
    to_signed(2, 8),
    to_signed(3, 8),
    to_signed(3, 8),
    to_signed(0, 8),
    to_signed(-4, 8),
    to_signed(-7, 8),
    to_signed(-10, 8),
    to_signed(-16, 8),
    to_signed(-24, 8),
    to_signed(-32, 8),
    to_signed(-40, 8),
    to_signed(-50, 8),
    to_signed(-61, 8),
    to_signed(-66, 8),
    to_signed(-60, 8),
    to_signed(-46, 8),
    to_signed(-30, 8),
    to_signed(-19, 8),
    to_signed(-13, 8),
    to_signed(-11, 8),
    to_signed(-7, 8),
    to_signed(-3, 8),
    to_signed(1, 8),
    to_signed(4, 8),
    to_signed(4, 8),
    to_signed(6, 8),
    to_signed(14, 8),
    to_signed(25, 8),
    to_signed(39, 8),
    to_signed(50, 8),
    to_signed(57, 8),
    to_signed(58, 8),
    to_signed(53, 8),
    to_signed(48, 8),
    to_signed(48, 8),
    to_signed(50, 8),
    to_signed(50, 8),
    to_signed(46, 8),
    to_signed(43, 8),
    to_signed(46, 8),
    to_signed(50, 8),
    to_signed(50, 8),
    to_signed(42, 8),
    to_signed(32, 8),
    to_signed(21, 8),
    to_signed(9, 8),
    to_signed(-3, 8),
    to_signed(-12, 8),
    to_signed(-14, 8),
    to_signed(-10, 8),
    to_signed(-5, 8),
    to_signed(-4, 8),
    to_signed(-7, 8),
    to_signed(-10, 8),
    to_signed(-11, 8),
    to_signed(-10, 8),
    to_signed(-9, 8),
    to_signed(-10, 8),
    to_signed(-12, 8),
    to_signed(-14, 8),
    to_signed(-13, 8),
    to_signed(-10, 8),
    to_signed(-6, 8),
    to_signed(1, 8),
    to_signed(10, 8),
    to_signed(20, 8),
    to_signed(29, 8),
    to_signed(36, 8),
    to_signed(38, 8),
    to_signed(34, 8),
    to_signed(26, 8),
    to_signed(16, 8),
    to_signed(4, 8),
    to_signed(-6, 8),
    to_signed(-12, 8),
    to_signed(-13, 8),
    to_signed(-12, 8),
    to_signed(-11, 8),
    to_signed(-10, 8),
    to_signed(-12, 8),
    to_signed(-17, 8),
    to_signed(-25, 8),
    to_signed(-36, 8),
    to_signed(-50, 8),
    to_signed(-66, 8),
    to_signed(-78, 8),
    to_signed(-83, 8),
    to_signed(-77, 8),
    to_signed(-65, 8),
    to_signed(-51, 8),
    to_signed(-38, 8),
    to_signed(-27, 8),
    to_signed(-19, 8),
    to_signed(-13, 8),
    to_signed(-9, 8),
    to_signed(-6, 8),
    to_signed(-4, 8),
    to_signed(1, 8),
    to_signed(10, 8),
    to_signed(21, 8),
    to_signed(32, 8),
    to_signed(46, 8),
    to_signed(60, 8),
    to_signed(73, 8),
    to_signed(78, 8),
    to_signed(75, 8),
    to_signed(70, 8),
    to_signed(69, 8),
    to_signed(73, 8),
    to_signed(76, 8),
    to_signed(74, 8),
    to_signed(65, 8),
    to_signed(56, 8),
    to_signed(47, 8),
    to_signed(40, 8),
    to_signed(29, 8),
    to_signed(14, 8),
    to_signed(-1, 8),
    to_signed(-12, 8),
    to_signed(-20, 8),
    to_signed(-25, 8),
    to_signed(-28, 8),
    to_signed(-29, 8),
    to_signed(-33, 8),
    to_signed(-41, 8),
    to_signed(-50, 8),
    to_signed(-51, 8),
    to_signed(-42, 8),
    to_signed(-30, 8),
    to_signed(-24, 8),
    to_signed(-26, 8),
    to_signed(-31, 8),
    to_signed(-31, 8),
    to_signed(-23, 8),
    to_signed(-7, 8),
    to_signed(10, 8),
    to_signed(22, 8),
    to_signed(30, 8),
    to_signed(34, 8),
    to_signed(35, 8),
    to_signed(31, 8),
    to_signed(21, 8),
    to_signed(10, 8),
    to_signed(1, 8),
    to_signed(-6, 8),
    to_signed(-10, 8),
    to_signed(-11, 8),
    to_signed(-9, 8),
    to_signed(-5, 8),
    to_signed(-3, 8),
    to_signed(-7, 8),
    to_signed(-20, 8),
    to_signed(-41, 8),
    to_signed(-63, 8),
    to_signed(-78, 8),
    to_signed(-83, 8),
    to_signed(-80, 8),
    to_signed(-74, 8),
    to_signed(-67, 8),
    to_signed(-60, 8),
    to_signed(-53, 8),
    to_signed(-45, 8),
    to_signed(-35, 8),
    to_signed(-25, 8),
    to_signed(-19, 8),
    to_signed(-18, 8),
    to_signed(-18, 8),
    to_signed(-14, 8),
    to_signed(-1, 8),
    to_signed(20, 8),
    to_signed(43, 8),
    to_signed(62, 8),
    to_signed(74, 8),
    to_signed(79, 8),
    to_signed(79, 8),
    to_signed(76, 8),
    to_signed(71, 8),
    to_signed(65, 8),
    to_signed(60, 8),
    to_signed(56, 8),
    to_signed(54, 8),
    to_signed(54, 8),
    to_signed(57, 8),
    to_signed(60, 8),
    to_signed(60, 8),
    to_signed(57, 8),
    to_signed(46, 8),
    to_signed(26, 8),
    to_signed(-1, 8),
    to_signed(-30, 8),
    to_signed(-51, 8),
    to_signed(-60, 8),
    to_signed(-57, 8),
    to_signed(-47, 8),
    to_signed(-37, 8),
    to_signed(-33, 8),
    to_signed(-36, 8),
    to_signed(-40, 8),
    to_signed(-39, 8),
    to_signed(-34, 8),
    to_signed(-32, 8),
    to_signed(-35, 8),
    to_signed(-40, 8),
    to_signed(-42, 8),
    to_signed(-41, 8),
    to_signed(-36, 8),
    to_signed(-23, 8),
    to_signed(-4, 8),
    to_signed(17, 8),
    to_signed(31, 8),
    to_signed(34, 8),
    to_signed(31, 8),
    to_signed(26, 8),
    to_signed(18, 8),
    to_signed(5, 8),
    to_signed(-10, 8),
    to_signed(-23, 8),
    to_signed(-29, 8),
    to_signed(-29, 8),
    to_signed(-26, 8),
    to_signed(-21, 8),
    to_signed(-14, 8),
    to_signed(-9, 8),
    to_signed(-12, 8),
    to_signed(-29, 8),
    to_signed(-54, 8),
    to_signed(-76, 8),
    to_signed(-87, 8),
    to_signed(-88, 8),
    to_signed(-85, 8),
    to_signed(-77, 8),
    to_signed(-66, 8),
    to_signed(-51, 8),
    to_signed(-37, 8),
    to_signed(-24, 8),
    to_signed(-13, 8),
    to_signed(-7, 8),
    to_signed(-5, 8),
    to_signed(-10, 8),
    to_signed(-15, 8),
    to_signed(-13, 8),
    to_signed(-1, 8),
    to_signed(20, 8),
    to_signed(43, 8),
    to_signed(60, 8),
    to_signed(73, 8),
    to_signed(80, 8),
    to_signed(81, 8),
    to_signed(72, 8),
    to_signed(56, 8),
    to_signed(41, 8),
    to_signed(33, 8),
    to_signed(31, 8),
    to_signed(29, 8),
    to_signed(27, 8),
    to_signed(27, 8),
    to_signed(35, 8),
    to_signed(47, 8),
    to_signed(54, 8),
    to_signed(52, 8),
    to_signed(41, 8),
    to_signed(23, 8),
    to_signed(4, 8),
    to_signed(-16, 8),
    to_signed(-34, 8),
    to_signed(-48, 8),
    to_signed(-53, 8),
    to_signed(-45, 8),
    to_signed(-27, 8),
    to_signed(-6, 8),
    to_signed(11, 8),
    to_signed(18, 8),
    to_signed(16, 8),
    to_signed(8, 8),
    to_signed(-2, 8),
    to_signed(-12, 8),
    to_signed(-22, 8),
    to_signed(-29, 8),
    to_signed(-30, 8),
    to_signed(-25, 8),
    to_signed(-14, 8),
    to_signed(2, 8),
    to_signed(16, 8),
    to_signed(24, 8),
    to_signed(24, 8),
    to_signed(17, 8),
    to_signed(11, 8),
    to_signed(7, 8),
    to_signed(1, 8),
    to_signed(-7, 8),
    to_signed(-17, 8),
    to_signed(-24, 8),
    to_signed(-26, 8),
    to_signed(-25, 8),
    to_signed(-22, 8),
    to_signed(-16, 8),
    to_signed(-8, 8),
    to_signed(-3, 8),
    to_signed(-5, 8),
    to_signed(-14, 8),
    to_signed(-26, 8),
    to_signed(-36, 8),
    to_signed(-46, 8),
    to_signed(-56, 8),
    to_signed(-63, 8),
    to_signed(-62, 8),
    to_signed(-49, 8),
    to_signed(-31, 8),
    to_signed(-15, 8),
    to_signed(-3, 8),
    to_signed(7, 8),
    to_signed(13, 8),
    to_signed(13, 8),
    to_signed(7, 8),
    to_signed(1, 8),
    to_signed(0, 8),
    to_signed(4, 8),
    to_signed(12, 8),
    to_signed(25, 8),
    to_signed(43, 8),
    to_signed(62, 8),
    to_signed(72, 8),
    to_signed(71, 8),
    to_signed(62, 8),
    to_signed(54, 8),
    to_signed(50, 8),
    to_signed(47, 8),
    to_signed(44, 8),
    to_signed(42, 8),
    to_signed(42, 8),
    to_signed(46, 8),
    to_signed(49, 8),
    to_signed(51, 8),
    to_signed(49, 8),
    to_signed(45, 8),
    to_signed(36, 8),
    to_signed(23, 8),
    to_signed(6, 8),
    to_signed(-13, 8),
    to_signed(-29, 8),
    to_signed(-38, 8),
    to_signed(-36, 8),
    to_signed(-27, 8),
    to_signed(-16, 8),
    to_signed(-7, 8),
    to_signed(-1, 8),
    to_signed(1, 8),
    to_signed(-1, 8),
    to_signed(-9, 8),
    to_signed(-23, 8),
    to_signed(-36, 8),
    to_signed(-43, 8),
    to_signed(-40, 8),
    to_signed(-31, 8),
    to_signed(-19, 8),
    to_signed(-6, 8),
    to_signed(6, 8),
    to_signed(15, 8),
    to_signed(17, 8),
    to_signed(14, 8),
    to_signed(8, 8),
    to_signed(3, 8),
    to_signed(-2, 8),
    to_signed(-8, 8),
    to_signed(-16, 8),
    to_signed(-23, 8),
    to_signed(-28, 8),
    to_signed(-30, 8),
    to_signed(-31, 8),
    to_signed(-30, 8),
    to_signed(-27, 8),
    to_signed(-26, 8),
    to_signed(-31, 8),
    to_signed(-41, 8),
    to_signed(-54, 8),
    to_signed(-65, 8),
    to_signed(-74, 8),
    to_signed(-83, 8),
    to_signed(-89, 8),
    to_signed(-89, 8),
    to_signed(-82, 8),
    to_signed(-69, 8),
    to_signed(-54, 8),
    to_signed(-41, 8),
    to_signed(-31, 8),
    to_signed(-25, 8),
    to_signed(-25, 8),
    to_signed(-28, 8),
    to_signed(-29, 8),
    to_signed(-21, 8),
    to_signed(-5, 8),
    to_signed(13, 8),
    to_signed(26, 8),
    to_signed(35, 8),
    to_signed(45, 8),
    to_signed(56, 8),
    to_signed(63, 8),
    to_signed(62, 8),
    to_signed(54, 8),
    to_signed(45, 8),
    to_signed(41, 8),
    to_signed(43, 8),
    to_signed(49, 8),
    to_signed(57, 8),
    to_signed(62, 8),
    to_signed(61, 8),
    to_signed(56, 8),
    to_signed(47, 8),
    to_signed(36, 8),
    to_signed(23, 8),
    to_signed(5, 8),
    to_signed(-16, 8),
    to_signed(-35, 8),
    to_signed(-46, 8),
    to_signed(-48, 8),
    to_signed(-41, 8),
    to_signed(-28, 8),
    to_signed(-14, 8),
    to_signed(-4, 8),
    to_signed(-1, 8),
    to_signed(-5, 8),
    to_signed(-14, 8),
    to_signed(-24, 8),
    to_signed(-32, 8),
    to_signed(-33, 8),
    to_signed(-27, 8),
    to_signed(-14, 8),
    to_signed(1, 8),
    to_signed(14, 8),
    to_signed(26, 8),
    to_signed(35, 8),
    to_signed(42, 8),
    to_signed(44, 8),
    to_signed(41, 8),
    to_signed(36, 8),
    to_signed(28, 8),
    to_signed(20, 8),
    to_signed(9, 8),
    to_signed(-2, 8),
    to_signed(-11, 8),
    to_signed(-15, 8),
    to_signed(-15, 8),
    to_signed(-12, 8),
    to_signed(-10, 8),
    to_signed(-9, 8),
    to_signed(-15, 8),
    to_signed(-27, 8),
    to_signed(-43, 8),
    to_signed(-57, 8),
    to_signed(-67, 8),
    to_signed(-73, 8),
    to_signed(-77, 8),
    to_signed(-76, 8),
    to_signed(-69, 8),
    to_signed(-58, 8),
    to_signed(-45, 8),
    to_signed(-33, 8),
    to_signed(-22, 8),
    to_signed(-10, 8),
    to_signed(-1, 8),
    to_signed(6, 8),
    to_signed(11, 8),
    to_signed(15, 8),
    to_signed(20, 8),
    to_signed(23, 8),
    to_signed(27, 8),
    to_signed(36, 8),
    to_signed(49, 8),
    to_signed(64, 8),
    to_signed(75, 8),
    to_signed(77, 8),
    to_signed(70, 8),
    to_signed(58, 8),
    to_signed(46, 8),
    to_signed(40, 8),
    to_signed(37, 8),
    to_signed(37, 8),
    to_signed(37, 8),
    to_signed(38, 8),
    to_signed(41, 8),
    to_signed(42, 8),
    to_signed(38, 8),
    to_signed(26, 8),
    to_signed(6, 8),
    to_signed(-18, 8),
    to_signed(-41, 8),
    to_signed(-58, 8),
    to_signed(-65, 8),
    to_signed(-61, 8),
    to_signed(-48, 8),
    to_signed(-31, 8),
    to_signed(-16, 8),
    to_signed(-8, 8),
    to_signed(-8, 8),
    to_signed(-13, 8),
    to_signed(-20, 8),
    to_signed(-26, 8),
    to_signed(-29, 8),
    to_signed(-27, 8),
    to_signed(-24, 8),
    to_signed(-20, 8),
    to_signed(-15, 8),
    to_signed(-6, 8),
    to_signed(6, 8),
    to_signed(18, 8),
    to_signed(24, 8),
    to_signed(24, 8),
    to_signed(20, 8),
    to_signed(16, 8),
    to_signed(11, 8),
    to_signed(4, 8),
    to_signed(-5, 8),
    to_signed(-15, 8),
    to_signed(-23, 8),
    to_signed(-29, 8),
    to_signed(-32, 8),
    to_signed(-31, 8),
    to_signed(-27, 8),
    to_signed(-24, 8),
    to_signed(-24, 8),
    to_signed(-28, 8),
    to_signed(-36, 8),
    to_signed(-47, 8),
    to_signed(-57, 8),
    to_signed(-64, 8),
    to_signed(-67, 8),
    to_signed(-65, 8),
    to_signed(-58, 8),
    to_signed(-47, 8),
    to_signed(-32, 8),
    to_signed(-14, 8),
    to_signed(6, 8),
    to_signed(21, 8),
    to_signed(29, 8),
    to_signed(29, 8),
    to_signed(25, 8),
    to_signed(24, 8),
    to_signed(31, 8),
    to_signed(43, 8),
    to_signed(55, 8),
    to_signed(65, 8),
    to_signed(73, 8),
    to_signed(81, 8),
    to_signed(86, 8),
    to_signed(87, 8),
    to_signed(82, 8),
    to_signed(74, 8),
    to_signed(66, 8),
    to_signed(59, 8),
    to_signed(56, 8),
    to_signed(54, 8),
    to_signed(54, 8),
    to_signed(52, 8),
    to_signed(45, 8),
    to_signed(32, 8),
    to_signed(14, 8),
    to_signed(-7, 8),
    to_signed(-26, 8),
    to_signed(-41, 8),
    to_signed(-51, 8),
    to_signed(-56, 8),
    to_signed(-55, 8),
    to_signed(-46, 8),
    to_signed(-34, 8),
    to_signed(-24, 8),
    to_signed(-23, 8),
    to_signed(-30, 8),
    to_signed(-39, 8),
    to_signed(-43, 8),
    to_signed(-41, 8),
    to_signed(-33, 8),
    to_signed(-25, 8),
    to_signed(-18, 8),
    to_signed(-12, 8),
    to_signed(-4, 8),
    to_signed(4, 8),
    to_signed(15, 8),
    to_signed(25, 8),
    to_signed(32, 8),
    to_signed(30, 8),
    to_signed(23, 8),
    to_signed(16, 8),
    to_signed(12, 8),
    to_signed(9, 8),
    to_signed(2, 8),
    to_signed(-11, 8),
    to_signed(-23, 8),
    to_signed(-31, 8),
    to_signed(-33, 8),
    to_signed(-34, 8),
    to_signed(-35, 8),
    to_signed(-37, 8),
    to_signed(-41, 8),
    to_signed(-46, 8),
    to_signed(-54, 8),
    to_signed(-65, 8),
    to_signed(-76, 8),
    to_signed(-86, 8),
    to_signed(-92, 8),
    to_signed(-94, 8),
    to_signed(-88, 8),
    to_signed(-74, 8),
    to_signed(-53, 8),
    to_signed(-28, 8),
    to_signed(-5, 8),
    to_signed(12, 8),
    to_signed(20, 8),
    to_signed(22, 8),
    to_signed(24, 8),
    to_signed(29, 8),
    to_signed(37, 8),
    to_signed(44, 8),
    to_signed(51, 8),
    to_signed(61, 8),
    to_signed(74, 8),
    to_signed(86, 8),
    to_signed(92, 8),
    to_signed(90, 8),
    to_signed(84, 8),
    to_signed(77, 8),
    to_signed(74, 8),
    to_signed(72, 8),
    to_signed(73, 8),
    to_signed(72, 8),
    to_signed(66, 8),
    to_signed(55, 8),
    to_signed(38, 8),
    to_signed(16, 8),
    to_signed(-8, 8),
    to_signed(-30, 8),
    to_signed(-46, 8),
    to_signed(-53, 8),
    to_signed(-50, 8),
    to_signed(-39, 8),
    to_signed(-26, 8),
    to_signed(-16, 8),
    to_signed(-14, 8),
    to_signed(-19, 8),
    to_signed(-29, 8),
    to_signed(-36, 8),
    to_signed(-37, 8),
    to_signed(-31, 8),
    to_signed(-22, 8),
    to_signed(-12, 8),
    to_signed(-2, 8),
    to_signed(11, 8),
    to_signed(27, 8),
    to_signed(41, 8),
    to_signed(50, 8),
    to_signed(52, 8),
    to_signed(50, 8),
    to_signed(46, 8),
    to_signed(42, 8),
    to_signed(36, 8),
    to_signed(30, 8),
    to_signed(21, 8),
    to_signed(12, 8),
    to_signed(4, 8),
    to_signed(-2, 8),
    to_signed(-4, 8),
    to_signed(-1, 8),
    to_signed(3, 8),
    to_signed(4, 8),
    to_signed(-3, 8),
    to_signed(-19, 8),
    to_signed(-40, 8),
    to_signed(-60, 8),
    to_signed(-73, 8),
    to_signed(-79, 8),
    to_signed(-75, 8),
    to_signed(-64, 8),
    to_signed(-51, 8),
    to_signed(-37, 8),
    to_signed(-25, 8),
    to_signed(-14, 8),
    to_signed(-4, 8),
    to_signed(3, 8),
    to_signed(6, 8),
    to_signed(5, 8),
    to_signed(5, 8),
    to_signed(10, 8),
    to_signed(22, 8),
    to_signed(40, 8),
    to_signed(58, 8),
    to_signed(72, 8),
    to_signed(81, 8),
    to_signed(83, 8),
    to_signed(79, 8),
    to_signed(71, 8),
    to_signed(64, 8),
    to_signed(61, 8),
    to_signed(60, 8),
    to_signed(59, 8),
    to_signed(55, 8),
    to_signed(50, 8),
    to_signed(46, 8),
    to_signed(43, 8),
    to_signed(40, 8),
    to_signed(32, 8),
    to_signed(13, 8),
    to_signed(-15, 8),
    to_signed(-42, 8),
    to_signed(-60, 8),
    to_signed(-63, 8),
    to_signed(-57, 8),
    to_signed(-45, 8),
    to_signed(-35, 8),
    to_signed(-28, 8),
    to_signed(-24, 8),
    to_signed(-21, 8),
    to_signed(-18, 8),
    to_signed(-17, 8),
    to_signed(-21, 8),
    to_signed(-26, 8),
    to_signed(-30, 8),
    to_signed(-26, 8),
    to_signed(-11, 8),
    to_signed(13, 8),
    to_signed(39, 8),
    to_signed(59, 8),
    to_signed(68, 8),
    to_signed(66, 8),
    to_signed(55, 8),
    to_signed(41, 8),
    to_signed(27, 8),
    to_signed(15, 8),
    to_signed(2, 8),
    to_signed(-11, 8),
    to_signed(-20, 8),
    to_signed(-21, 8),
    to_signed(-13, 8),
    to_signed(-2, 8),
    to_signed(5, 8),
    to_signed(5, 8),
    to_signed(-4, 8),
    to_signed(-20, 8),
    to_signed(-42, 8),
    to_signed(-65, 8),
    to_signed(-81, 8),
    to_signed(-86, 8),
    to_signed(-82, 8),
    to_signed(-71, 8),
    to_signed(-59, 8),
    to_signed(-45, 8),
    to_signed(-31, 8),
    to_signed(-20, 8),
    to_signed(-14, 8),
    to_signed(-13, 8),
    to_signed(-12, 8),
    to_signed(-8, 8),
    to_signed(-1, 8),
    to_signed(6, 8),
    to_signed(13, 8),
    to_signed(23, 8),
    to_signed(36, 8),
    to_signed(52, 8),
    to_signed(64, 8),
    to_signed(68, 8),
    to_signed(64, 8),
    to_signed(55, 8),
    to_signed(43, 8),
    to_signed(32, 8),
    to_signed(25, 8),
    to_signed(20, 8),
    to_signed(19, 8),
    to_signed(19, 8),
    to_signed(20, 8),
    to_signed(21, 8),
    to_signed(20, 8),
    to_signed(17, 8),
    to_signed(10, 8),
    to_signed(-3, 8),
    to_signed(-24, 8),
    to_signed(-48, 8),
    to_signed(-69, 8),
    to_signed(-78, 8),
    to_signed(-74, 8),
    to_signed(-58, 8),
    to_signed(-37, 8),
    to_signed(-18, 8),
    to_signed(-8, 8),
    to_signed(-7, 8),
    to_signed(-9, 8),
    to_signed(-11, 8),
    to_signed(-12, 8),
    to_signed(-13, 8),
    to_signed(-17, 8),
    to_signed(-21, 8),
    to_signed(-19, 8),
    to_signed(-6, 8),
    to_signed(16, 8),
    to_signed(38, 8),
    to_signed(51, 8),
    to_signed(51, 8),
    to_signed(43, 8),
    to_signed(28, 8),
    to_signed(12, 8),
    to_signed(-4, 8),
    to_signed(-19, 8),
    to_signed(-33, 8),
    to_signed(-44, 8),
    to_signed(-50, 8),
    to_signed(-48, 8),
    to_signed(-42, 8),
    to_signed(-34, 8),
    to_signed(-27, 8),
    to_signed(-24, 8),
    to_signed(-28, 8),
    to_signed(-39, 8),
    to_signed(-57, 8),
    to_signed(-77, 8),
    to_signed(-92, 8),
    to_signed(-95, 8),
    to_signed(-86, 8),
    to_signed(-70, 8),
    to_signed(-51, 8),
    to_signed(-35, 8),
    to_signed(-20, 8),
    to_signed(-6, 8),
    to_signed(5, 8),
    to_signed(11, 8),
    to_signed(12, 8),
    to_signed(10, 8),
    to_signed(6, 8),
    to_signed(2, 8),
    to_signed(2, 8),
    to_signed(9, 8),
    to_signed(22, 8),
    to_signed(36, 8),
    to_signed(47, 8),
    to_signed(50, 8),
    to_signed(47, 8),
    to_signed(39, 8),
    to_signed(27, 8),
    to_signed(17, 8),
    to_signed(8, 8),
    to_signed(1, 8),
    to_signed(-4, 8),
    to_signed(-7, 8),
    to_signed(-8, 8),
    to_signed(-6, 8),
    to_signed(1, 8),
    to_signed(12, 8),
    to_signed(21, 8),
    to_signed(21, 8),
    to_signed(9, 8),
    to_signed(-9, 8),
    to_signed(-24, 8),
    to_signed(-32, 8),
    to_signed(-32, 8),
    to_signed(-27, 8),
    to_signed(-20, 8),
    to_signed(-9, 8),
    to_signed(4, 8),
    to_signed(18, 8),
    to_signed(30, 8),
    to_signed(36, 8),
    to_signed(34, 8),
    to_signed(25, 8),
    to_signed(10, 8),
    to_signed(-3, 8),
    to_signed(-9, 8),
    to_signed(-5, 8),
    to_signed(6, 8),
    to_signed(17, 8),
    to_signed(26, 8),
    to_signed(31, 8),
    to_signed(30, 8),
    to_signed(22, 8),
    to_signed(9, 8),
    to_signed(-6, 8),
    to_signed(-18, 8),
    to_signed(-28, 8),
    to_signed(-35, 8),
    to_signed(-38, 8),
    to_signed(-36, 8),
    to_signed(-29, 8),
    to_signed(-19, 8),
    to_signed(-9, 8),
    to_signed(-4, 8),
    to_signed(-3, 8),
    to_signed(-8, 8),
    to_signed(-17, 8),
    to_signed(-29, 8),
    to_signed(-39, 8),
    to_signed(-41, 8),
    to_signed(-34, 8),
    to_signed(-25, 8),
    to_signed(-17, 8),
    to_signed(-11, 8),
    to_signed(-4, 8),
    to_signed(5, 8),
    to_signed(16, 8),
    to_signed(26, 8),
    to_signed(32, 8),
    to_signed(30, 8),
    to_signed(23, 8),
    to_signed(16, 8),
    to_signed(15, 8),
    to_signed(19, 8),
    to_signed(27, 8),
    to_signed(37, 8),
    to_signed(48, 8),
    to_signed(56, 8),
    to_signed(62, 8),
    to_signed(66, 8),
    to_signed(68, 8),
    to_signed(68, 8),
    to_signed(63, 8),
    to_signed(53, 8),
    to_signed(42, 8),
    to_signed(35, 8),
    to_signed(35, 8),
    to_signed(41, 8),
    to_signed(52, 8),
    to_signed(63, 8),
    to_signed(70, 8),
    to_signed(67, 8),
    to_signed(54, 8),
    to_signed(34, 8),
    to_signed(14, 8),
    to_signed(-3, 8),
    to_signed(-17, 8),
    to_signed(-27, 8),
    to_signed(-31, 8),
    to_signed(-27, 8),
    to_signed(-14, 8),
    to_signed(5, 8),
    to_signed(23, 8),
    to_signed(33, 8),
    to_signed(32, 8),
    to_signed(20, 8),
    to_signed(1, 8),
    to_signed(-16, 8),
    to_signed(-25, 8),
    to_signed(-24, 8),
    to_signed(-16, 8),
    to_signed(-3, 8),
    to_signed(9, 8),
    to_signed(20, 8),
    to_signed(29, 8),
    to_signed(35, 8),
    to_signed(35, 8),
    to_signed(28, 8),
    to_signed(14, 8),
    to_signed(-3, 8),
    to_signed(-17, 8),
    to_signed(-23, 8),
    to_signed(-22, 8),
    to_signed(-18, 8),
    to_signed(-15, 8),
    to_signed(-15, 8),
    to_signed(-19, 8),
    to_signed(-26, 8),
    to_signed(-34, 8),
    to_signed(-43, 8),
    to_signed(-48, 8),
    to_signed(-50, 8),
    to_signed(-51, 8),
    to_signed(-56, 8),
    to_signed(-65, 8),
    to_signed(-70, 8),
    to_signed(-67, 8),
    to_signed(-56, 8),
    to_signed(-43, 8),
    to_signed(-31, 8),
    to_signed(-20, 8),
    to_signed(-9, 8),
    to_signed(3, 8),
    to_signed(16, 8),
    to_signed(29, 8),
    to_signed(40, 8),
    to_signed(46, 8),
    to_signed(47, 8),
    to_signed(49, 8),
    to_signed(55, 8),
    to_signed(64, 8),
    to_signed(71, 8),
    to_signed(75, 8),
    to_signed(75, 8),
    to_signed(72, 8),
    to_signed(66, 8),
    to_signed(60, 8),
    to_signed(55, 8),
    to_signed(50, 8),
    to_signed(47, 8),
    to_signed(45, 8),
    to_signed(43, 8),
    to_signed(39, 8),
    to_signed(31, 8),
    to_signed(17, 8),
    to_signed(0, 8),
    to_signed(-20, 8),
    to_signed(-40, 8),
    to_signed(-60, 8),
    to_signed(-75, 8),
    to_signed(-79, 8),
    to_signed(-70, 8),
    to_signed(-53, 8),
    to_signed(-35, 8),
    to_signed(-21, 8),
    to_signed(-14, 8),
    to_signed(-11, 8),
    to_signed(-14, 8),
    to_signed(-21, 8),
    to_signed(-30, 8),
    to_signed(-34, 8),
    to_signed(-31, 8),
    to_signed(-22, 8),
    to_signed(-11, 8),
    to_signed(1, 8),
    to_signed(13, 8),
    to_signed(24, 8),
    to_signed(28, 8),
    to_signed(24, 8),
    to_signed(15, 8),
    to_signed(4, 8),
    to_signed(-7, 8),
    to_signed(-19, 8),
    to_signed(-30, 8),
    to_signed(-39, 8),
    to_signed(-46, 8),
    to_signed(-51, 8),
    to_signed(-56, 8),
    to_signed(-60, 8),
    to_signed(-63, 8),
    to_signed(-67, 8),
    to_signed(-75, 8),
    to_signed(-84, 8),
    to_signed(-93, 8),
    to_signed(-97, 8),
    to_signed(-97, 8),
    to_signed(-95, 8),
    to_signed(-92, 8),
    to_signed(-85, 8),
    to_signed(-72, 8),
    to_signed(-56, 8),
    to_signed(-37, 8),
    to_signed(-17, 8),
    to_signed(0, 8),
    to_signed(14, 8),
    to_signed(24, 8),
    to_signed(36, 8),
    to_signed(50, 8),
    to_signed(63, 8),
    to_signed(70, 8),
    to_signed(72, 8),
    to_signed(72, 8),
    to_signed(73, 8),
    to_signed(75, 8),
    to_signed(78, 8),
    to_signed(79, 8),
    to_signed(76, 8),
    to_signed(69, 8),
    to_signed(59, 8),
    to_signed(51, 8),
    to_signed(47, 8),
    to_signed(44, 8),
    to_signed(42, 8),
    to_signed(39, 8),
    to_signed(35, 8),
    to_signed(30, 8),
    to_signed(23, 8),
    to_signed(11, 8),
    to_signed(-8, 8),
    to_signed(-30, 8),
    to_signed(-50, 8),
    to_signed(-62, 8),
    to_signed(-65, 8),
    to_signed(-60, 8),
    to_signed(-47, 8),
    to_signed(-31, 8),
    to_signed(-13, 8),
    to_signed(2, 8),
    to_signed(10, 8),
    to_signed(11, 8),
    to_signed(5, 8),
    to_signed(-3, 8),
    to_signed(-9, 8),
    to_signed(-11, 8),
    to_signed(-10, 8),
    to_signed(-7, 8),
    to_signed(-1, 8),
    to_signed(10, 8),
    to_signed(26, 8),
    to_signed(38, 8),
    to_signed(41, 8),
    to_signed(33, 8),
    to_signed(18, 8),
    to_signed(2, 8),
    to_signed(-11, 8),
    to_signed(-22, 8),
    to_signed(-30, 8),
    to_signed(-37, 8),
    to_signed(-42, 8),
    to_signed(-46, 8),
    to_signed(-48, 8),
    to_signed(-48, 8),
    to_signed(-49, 8),
    to_signed(-53, 8),
    to_signed(-60, 8),
    to_signed(-68, 8),
    to_signed(-72, 8),
    to_signed(-71, 8),
    to_signed(-67, 8),
    to_signed(-63, 8),
    to_signed(-59, 8),
    to_signed(-53, 8),
    to_signed(-46, 8),
    to_signed(-37, 8),
    to_signed(-25, 8),
    to_signed(-10, 8),
    to_signed(7, 8),
    to_signed(25, 8),
    to_signed(39, 8),
    to_signed(49, 8),
    to_signed(54, 8),
    to_signed(53, 8),
    to_signed(49, 8),
    to_signed(45, 8),
    to_signed(43, 8),
    to_signed(42, 8),
    to_signed(42, 8),
    to_signed(43, 8),
    to_signed(45, 8),
    to_signed(48, 8),
    to_signed(53, 8),
    to_signed(58, 8),
    to_signed(60, 8),
    to_signed(56, 8),
    to_signed(47, 8),
    to_signed(37, 8),
    to_signed(27, 8),
    to_signed(18, 8),
    to_signed(6, 8),
    to_signed(-8, 8),
    to_signed(-23, 8),
    to_signed(-38, 8),
    to_signed(-50, 8),
    to_signed(-57, 8),
    to_signed(-56, 8),
    to_signed(-50, 8),
    to_signed(-39, 8),
    to_signed(-28, 8),
    to_signed(-20, 8),
    to_signed(-15, 8),
    to_signed(-14, 8),
    to_signed(-17, 8),
    to_signed(-21, 8),
    to_signed(-23, 8),
    to_signed(-21, 8),
    to_signed(-17, 8),
    to_signed(-12, 8),
    to_signed(-4, 8),
    to_signed(6, 8),
    to_signed(17, 8),
    to_signed(26, 8),
    to_signed(27, 8),
    to_signed(19, 8),
    to_signed(5, 8),
    to_signed(-8, 8),
    to_signed(-17, 8),
    to_signed(-21, 8),
    to_signed(-22, 8),
    to_signed(-23, 8),
    to_signed(-24, 8),
    to_signed(-25, 8),
    to_signed(-29, 8),
    to_signed(-35, 8),
    to_signed(-42, 8),
    to_signed(-47, 8),
    to_signed(-48, 8),
    to_signed(-47, 8),
    to_signed(-47, 8),
    to_signed(-48, 8),
    to_signed(-50, 8),
    to_signed(-48, 8),
    to_signed(-44, 8),
    to_signed(-38, 8),
    to_signed(-33, 8),
    to_signed(-27, 8),
    to_signed(-19, 8),
    to_signed(-7, 8),
    to_signed(6, 8),
    to_signed(19, 8),
    to_signed(30, 8),
    to_signed(39, 8),
    to_signed(45, 8),
    to_signed(49, 8),
    to_signed(52, 8),
    to_signed(56, 8),
    to_signed(60, 8),
    to_signed(61, 8),
    to_signed(59, 8),
    to_signed(56, 8),
    to_signed(53, 8),
    to_signed(48, 8),
    to_signed(43, 8),
    to_signed(40, 8),
    to_signed(43, 8),
    to_signed(51, 8),
    to_signed(58, 8),
    to_signed(58, 8),
    to_signed(50, 8),
    to_signed(37, 8),
    to_signed(20, 8),
    to_signed(-2, 8),
    to_signed(-27, 8),
    to_signed(-51, 8),
    to_signed(-68, 8),
    to_signed(-78, 8),
    to_signed(-78, 8),
    to_signed(-64, 8),
    to_signed(-42, 8),
    to_signed(-20, 8),
    to_signed(-7, 8),
    to_signed(-4, 8),
    to_signed(-9, 8),
    to_signed(-19, 8),
    to_signed(-30, 8),
    to_signed(-40, 8),
    to_signed(-42, 8),
    to_signed(-36, 8),
    to_signed(-22, 8),
    to_signed(-4, 8),
    to_signed(16, 8),
    to_signed(35, 8),
    to_signed(48, 8),
    to_signed(54, 8),
    to_signed(51, 8),
    to_signed(40, 8),
    to_signed(23, 8),
    to_signed(4, 8),
    to_signed(-12, 8),
    to_signed(-22, 8),
    to_signed(-26, 8),
    to_signed(-26, 8),
    to_signed(-24, 8),
    to_signed(-19, 8),
    to_signed(-12, 8),
    to_signed(-6, 8),
    to_signed(-7, 8),
    to_signed(-14, 8),
    to_signed(-27, 8),
    to_signed(-40, 8),
    to_signed(-51, 8),
    to_signed(-59, 8),
    to_signed(-61, 8),
    to_signed(-55, 8),
    to_signed(-42, 8),
    to_signed(-25, 8),
    to_signed(-9, 8),
    to_signed(5, 8),
    to_signed(17, 8),
    to_signed(27, 8),
    to_signed(33, 8),
    to_signed(35, 8),
    to_signed(36, 8),
    to_signed(41, 8),
    to_signed(50, 8),
    to_signed(59, 8),
    to_signed(66, 8),
    to_signed(71, 8),
    to_signed(77, 8),
    to_signed(81, 8),
    to_signed(78, 8),
    to_signed(68, 8),
    to_signed(54, 8),
    to_signed(40, 8),
    to_signed(31, 8),
    to_signed(27, 8),
    to_signed(29, 8),
    to_signed(35, 8),
    to_signed(41, 8),
    to_signed(44, 8),
    to_signed(43, 8),
    to_signed(38, 8),
    to_signed(29, 8),
    to_signed(11, 8),
    to_signed(-15, 8),
    to_signed(-41, 8),
    to_signed(-59, 8),
    to_signed(-63, 8),
    to_signed(-52, 8),
    to_signed(-31, 8),
    to_signed(-4, 8),
    to_signed(18, 8),
    to_signed(30, 8),
    to_signed(32, 8),
    to_signed(28, 8),
    to_signed(22, 8),
    to_signed(14, 8),
    to_signed(5, 8),
    to_signed(-1, 8),
    to_signed(0, 8),
    to_signed(9, 8),
    to_signed(26, 8),
    to_signed(48, 8),
    to_signed(66, 8),
    to_signed(73, 8),
    to_signed(69, 8),
    to_signed(55, 8),
    to_signed(37, 8),
    to_signed(20, 8),
    to_signed(5, 8),
    to_signed(-7, 8),
    to_signed(-17, 8),
    to_signed(-25, 8),
    to_signed(-30, 8),
    to_signed(-28, 8),
    to_signed(-21, 8),
    to_signed(-14, 8),
    to_signed(-12, 8),
    to_signed(-16, 8),
    to_signed(-26, 8),
    to_signed(-38, 8),
    to_signed(-50, 8),
    to_signed(-59, 8),
    to_signed(-61, 8),
    to_signed(-56, 8),
    to_signed(-47, 8),
    to_signed(-35, 8),
    to_signed(-23, 8),
    to_signed(-10, 8),
    to_signed(3, 8),
    to_signed(16, 8),
    to_signed(28, 8),
    to_signed(39, 8),
    to_signed(45, 8),
    to_signed(46, 8),
    to_signed(41, 8),
    to_signed(37, 8),
    to_signed(37, 8),
    to_signed(42, 8),
    to_signed(52, 8),
    to_signed(62, 8),
    to_signed(65, 8),
    to_signed(61, 8),
    to_signed(51, 8),
    to_signed(40, 8),
    to_signed(31, 8),
    to_signed(23, 8),
    to_signed(12, 8),
    to_signed(2, 8),
    to_signed(-4, 8),
    to_signed(-4, 8),
    to_signed(1, 8),
    to_signed(10, 8),
    to_signed(19, 8),
    to_signed(22, 8),
    to_signed(15, 8),
    to_signed(-4, 8),
    to_signed(-28, 8),
    to_signed(-49, 8),
    to_signed(-62, 8),
    to_signed(-64, 8),
    to_signed(-57, 8),
    to_signed(-44, 8),
    to_signed(-27, 8),
    to_signed(-9, 8),
    to_signed(10, 8),
    to_signed(24, 8),
    to_signed(30, 8),
    to_signed(26, 8),
    to_signed(14, 8),
    to_signed(-2, 8),
    to_signed(-18, 8),
    to_signed(-26, 8),
    to_signed(-20, 8),
    to_signed(-2, 8),
    to_signed(21, 8),
    to_signed(36, 8),
    to_signed(40, 8),
    to_signed(34, 8),
    to_signed(23, 8),
    to_signed(5, 8),
    to_signed(-18, 8),
    to_signed(-40, 8),
    to_signed(-57, 8),
    to_signed(-67, 8),
    to_signed(-72, 8),
    to_signed(-71, 8),
    to_signed(-63, 8),
    to_signed(-51, 8),
    to_signed(-40, 8),
    to_signed(-36, 8),
    to_signed(-41, 8),
    to_signed(-57, 8),
    to_signed(-76, 8),
    to_signed(-89, 8),
    to_signed(-93, 8),
    to_signed(-88, 8),
    to_signed(-81, 8),
    to_signed(-71, 8),
    to_signed(-58, 8),
    to_signed(-41, 8),
    to_signed(-22, 8),
    to_signed(-4, 8),
    to_signed(9, 8),
    to_signed(17, 8),
    to_signed(18, 8),
    to_signed(13, 8),
    to_signed(7, 8),
    to_signed(6, 8),
    to_signed(10, 8),
    to_signed(18, 8),
    to_signed(27, 8),
    to_signed(34, 8),
    to_signed(41, 8),
    to_signed(43, 8),
    to_signed(38, 8),
    to_signed(26, 8),
    to_signed(12, 8),
    to_signed(1, 8),
    to_signed(-8, 8),
    to_signed(-13, 8),
    to_signed(-16, 8),
    to_signed(-16, 8),
    to_signed(-12, 8),
    to_signed(-4, 8),
    to_signed(5, 8),
    to_signed(13, 8),
    to_signed(14, 8),
    to_signed(5, 8),
    to_signed(-12, 8),
    to_signed(-35, 8),
    to_signed(-56, 8),
    to_signed(-71, 8),
    to_signed(-76, 8),
    to_signed(-74, 8),
    to_signed(-67, 8),
    to_signed(-53, 8),
    to_signed(-36, 8),
    to_signed(-17, 8),
    to_signed(-3, 8),
    to_signed(5, 8),
    to_signed(7, 8),
    to_signed(2, 8),
    to_signed(-9, 8),
    to_signed(-24, 8),
    to_signed(-34, 8),
    to_signed(-34, 8),
    to_signed(-25, 8),
    to_signed(-15, 8),
    to_signed(-9, 8),
    to_signed(-6, 8),
    to_signed(-6, 8),
    to_signed(-9, 8),
    to_signed(-15, 8),
    to_signed(-23, 8),
    to_signed(-32, 8),
    to_signed(-43, 8),
    to_signed(-53, 8),
    to_signed(-59, 8),
    to_signed(-59, 8),
    to_signed(-53, 8),
    to_signed(-47, 8),
    to_signed(-42, 8),
    to_signed(-42, 8),
    to_signed(-48, 8),
    to_signed(-55, 8),
    to_signed(-59, 8),
    to_signed(-56, 8),
    to_signed(-50, 8),
    to_signed(-44, 8),
    to_signed(-39, 8),
    to_signed(-33, 8),
    to_signed(-27, 8),
    to_signed(-25, 8),
    to_signed(-25, 8),
    to_signed(-22, 8),
    to_signed(-15, 8),
    to_signed(-7, 8),
    to_signed(2, 8),
    to_signed(12, 8),
    to_signed(23, 8),
    to_signed(34, 8),
    to_signed(42, 8),
    to_signed(47, 8),
    to_signed(47, 8),
    to_signed(42, 8),
    to_signed(34, 8),
    to_signed(25, 8),
    to_signed(21, 8),
    to_signed(22, 8),
    to_signed(27, 8),
    to_signed(32, 8),
    to_signed(35, 8),
    to_signed(37, 8),
    to_signed(39, 8),
    to_signed(40, 8),
    to_signed(40, 8),
    to_signed(42, 8),
    to_signed(46, 8),
    to_signed(48, 8),
    to_signed(46, 8),
    to_signed(42, 8),
    to_signed(34, 8),
    to_signed(21, 8),
    to_signed(4, 8),
    to_signed(-13, 8),
    to_signed(-26, 8),
    to_signed(-34, 8),
    to_signed(-35, 8),
    to_signed(-29, 8),
    to_signed(-16, 8),
    to_signed(0, 8),
    to_signed(14, 8),
    to_signed(23, 8),
    to_signed(23, 8),
    to_signed(15, 8),
    to_signed(2, 8),
    to_signed(-9, 8),
    to_signed(-16, 8),
    to_signed(-16, 8),
    to_signed(-9, 8),
    to_signed(2, 8),
    to_signed(14, 8),
    to_signed(22, 8),
    to_signed(22, 8),
    to_signed(18, 8),
    to_signed(11, 8),
    to_signed(2, 8),
    to_signed(-8, 8),
    to_signed(-15, 8),
    to_signed(-17, 8),
    to_signed(-15, 8),
    to_signed(-15, 8),
    to_signed(-16, 8),
    to_signed(-15, 8),
    to_signed(-12, 8),
    to_signed(-13, 8),
    to_signed(-23, 8),
    to_signed(-33, 8),
    to_signed(-37, 8),
    to_signed(-34, 8),
    to_signed(-27, 8),
    to_signed(-20, 8),
    to_signed(-13, 8),
    to_signed(-9, 8),
    to_signed(-10, 8),
    to_signed(-14, 8),
    to_signed(-14, 8),
    to_signed(-9, 8),
    to_signed(-2, 8),
    to_signed(5, 8),
    to_signed(16, 8),
    to_signed(31, 8),
    to_signed(50, 8),
    to_signed(68, 8),
    to_signed(81, 8),
    to_signed(88, 8),
    to_signed(87, 8),
    to_signed(79, 8),
    to_signed(66, 8),
    to_signed(56, 8),
    to_signed(50, 8),
    to_signed(51, 8),
    to_signed(57, 8),
    to_signed(66, 8),
    to_signed(78, 8),
    to_signed(89, 8),
    to_signed(96, 8),
    to_signed(98, 8),
    to_signed(95, 8),
    to_signed(88, 8),
    to_signed(76, 8),
    to_signed(63, 8),
    to_signed(52, 8),
    to_signed(41, 8),
    to_signed(29, 8),
    to_signed(14, 8),
    to_signed(-4, 8),
    to_signed(-19, 8),
    to_signed(-27, 8),
    to_signed(-30, 8),
    to_signed(-27, 8),
    to_signed(-19, 8),
    to_signed(-9, 8),
    to_signed(-2, 8),
    to_signed(2, 8),
    to_signed(1, 8),
    to_signed(-2, 8),
    to_signed(-7, 8),
    to_signed(-13, 8),
    to_signed(-16, 8),
    to_signed(-10, 8),
    to_signed(3, 8),
    to_signed(18, 8),
    to_signed(30, 8),
    to_signed(34, 8),
    to_signed(31, 8),
    to_signed(24, 8),
    to_signed(16, 8),
    to_signed(5, 8),
    to_signed(-6, 8),
    to_signed(-14, 8),
    to_signed(-16, 8),
    to_signed(-12, 8),
    to_signed(-8, 8),
    to_signed(-6, 8),
    to_signed(-6, 8),
    to_signed(-9, 8),
    to_signed(-18, 8),
    to_signed(-33, 8),
    to_signed(-45, 8),
    to_signed(-50, 8),
    to_signed(-50, 8),
    to_signed(-47, 8),
    to_signed(-43, 8),
    to_signed(-36, 8),
    to_signed(-29, 8),
    to_signed(-27, 8),
    to_signed(-27, 8),
    to_signed(-25, 8),
    to_signed(-21, 8),
    to_signed(-16, 8),
    to_signed(-8, 8),
    to_signed(4, 8),
    to_signed(21, 8),
    to_signed(39, 8),
    to_signed(54, 8),
    to_signed(64, 8),
    to_signed(70, 8),
    to_signed(69, 8),
    to_signed(62, 8),
    to_signed(53, 8),
    to_signed(45, 8),
    to_signed(40, 8),
    to_signed(40, 8),
    to_signed(43, 8),
    to_signed(47, 8),
    to_signed(52, 8),
    to_signed(59, 8),
    to_signed(66, 8),
    to_signed(72, 8),
    to_signed(73, 8),
    to_signed(69, 8),
    to_signed(58, 8),
    to_signed(43, 8),
    to_signed(24, 8),
    to_signed(7, 8),
    to_signed(-11, 8),
    to_signed(-29, 8),
    to_signed(-50, 8),
    to_signed(-68, 8),
    to_signed(-76, 8),
    to_signed(-72, 8),
    to_signed(-56, 8),
    to_signed(-35, 8),
    to_signed(-15, 8),
    to_signed(-2, 8),
    to_signed(3, 8),
    to_signed(1, 8),
    to_signed(-5, 8),
    to_signed(-11, 8),
    to_signed(-15, 8),
    to_signed(-16, 8),
    to_signed(-12, 8),
    to_signed(-5, 8),
    to_signed(8, 8),
    to_signed(23, 8),
    to_signed(35, 8),
    to_signed(40, 8),
    to_signed(36, 8),
    to_signed(27, 8),
    to_signed(14, 8),
    to_signed(-2, 8),
    to_signed(-18, 8),
    to_signed(-29, 8),
    to_signed(-33, 8),
    to_signed(-32, 8),
    to_signed(-32, 8),
    to_signed(-33, 8),
    to_signed(-34, 8),
    to_signed(-37, 8),
    to_signed(-43, 8),
    to_signed(-48, 8),
    to_signed(-53, 8),
    to_signed(-56, 8),
    to_signed(-58, 8),
    to_signed(-59, 8),
    to_signed(-58, 8),
    to_signed(-57, 8),
    to_signed(-57, 8),
    to_signed(-55, 8),
    to_signed(-50, 8),
    to_signed(-42, 8),
    to_signed(-32, 8),
    to_signed(-18, 8),
    to_signed(1, 8),
    to_signed(20, 8),
    to_signed(33, 8),
    to_signed(40, 8),
    to_signed(44, 8),
    to_signed(46, 8),
    to_signed(47, 8),
    to_signed(46, 8),
    to_signed(45, 8),
    to_signed(43, 8),
    to_signed(41, 8),
    to_signed(40, 8),
    to_signed(40, 8),
    to_signed(43, 8),
    to_signed(48, 8),
    to_signed(52, 8),
    to_signed(57, 8),
    to_signed(60, 8),
    to_signed(61, 8),
    to_signed(57, 8),
    to_signed(48, 8),
    to_signed(31, 8),
    to_signed(7, 8),
    to_signed(-23, 8),
    to_signed(-52, 8),
    to_signed(-77, 8),
    to_signed(-94, 8),
    to_signed(-98, 8),
    to_signed(-88, 8),
    to_signed(-67, 8),
    to_signed(-41, 8),
    to_signed(-18, 8),
    to_signed(-1, 8),
    to_signed(6, 8),
    to_signed(3, 8),
    to_signed(-10, 8),
    to_signed(-26, 8),
    to_signed(-37, 8),
    to_signed(-38, 8),
    to_signed(-29, 8),
    to_signed(-13, 8),
    to_signed(8, 8),
    to_signed(29, 8),
    to_signed(44, 8),
    to_signed(51, 8),
    to_signed(48, 8),
    to_signed(38, 8),
    to_signed(23, 8),
    to_signed(5, 8),
    to_signed(-15, 8),
    to_signed(-35, 8),
    to_signed(-49, 8),
    to_signed(-54, 8),
    to_signed(-53, 8),
    to_signed(-49, 8),
    to_signed(-44, 8),
    to_signed(-38, 8),
    to_signed(-34, 8),
    to_signed(-35, 8),
    to_signed(-42, 8),
    to_signed(-50, 8),
    to_signed(-59, 8),
    to_signed(-67, 8),
    to_signed(-72, 8),
    to_signed(-73, 8),
    to_signed(-71, 8),
    to_signed(-65, 8),
    to_signed(-53, 8),
    to_signed(-35, 8),
    to_signed(-11, 8),
    to_signed(11, 8),
    to_signed(28, 8),
    to_signed(38, 8),
    to_signed(44, 8),
    to_signed(48, 8),
    to_signed(52, 8),
    to_signed(56, 8),
    to_signed(60, 8),
    to_signed(61, 8),
    to_signed(58, 8),
    to_signed(54, 8),
    to_signed(51, 8),
    to_signed(48, 8),
    to_signed(45, 8),
    to_signed(44, 8),
    to_signed(43, 8),
    to_signed(42, 8),
    to_signed(41, 8),
    to_signed(42, 8),
    to_signed(41, 8),
    to_signed(36, 8),
    to_signed(25, 8),
    to_signed(10, 8),
    to_signed(-8, 8),
    to_signed(-29, 8),
    to_signed(-52, 8),
    to_signed(-74, 8),
    to_signed(-89, 8),
    to_signed(-91, 8),
    to_signed(-80, 8),
    to_signed(-59, 8),
    to_signed(-33, 8),
    to_signed(-9, 8),
    to_signed(7, 8),
    to_signed(15, 8),
    to_signed(15, 8),
    to_signed(8, 8),
    to_signed(-4, 8),
    to_signed(-16, 8),
    to_signed(-22, 8),
    to_signed(-17, 8),
    to_signed(-2, 8),
    to_signed(22, 8),
    to_signed(48, 8),
    to_signed(66, 8),
    to_signed(73, 8),
    to_signed(67, 8),
    to_signed(52, 8),
    to_signed(33, 8),
    to_signed(12, 8),
    to_signed(-9, 8),
    to_signed(-28, 8),
    to_signed(-42, 8),
    to_signed(-50, 8),
    to_signed(-52, 8),
    to_signed(-47, 8),
    to_signed(-40, 8),
    to_signed(-33, 8),
    to_signed(-31, 8),
    to_signed(-33, 8),
    to_signed(-38, 8),
    to_signed(-45, 8),
    to_signed(-50, 8),
    to_signed(-54, 8),
    to_signed(-55, 8),
    to_signed(-53, 8),
    to_signed(-47, 8),
    to_signed(-38, 8),
    to_signed(-25, 8),
    to_signed(-9, 8),
    to_signed(12, 8),
    to_signed(33, 8),
    to_signed(48, 8),
    to_signed(55, 8),
    to_signed(58, 8),
    to_signed(60, 8),
    to_signed(63, 8),
    to_signed(64, 8),
    to_signed(66, 8),
    to_signed(68, 8),
    to_signed(69, 8),
    to_signed(68, 8),
    to_signed(60, 8),
    to_signed(50, 8),
    to_signed(40, 8),
    to_signed(31, 8),
    to_signed(25, 8),
    to_signed(20, 8),
    to_signed(18, 8),
    to_signed(19, 8),
    to_signed(22, 8),
    to_signed(24, 8),
    to_signed(23, 8),
    to_signed(21, 8),
    to_signed(17, 8),
    to_signed(7, 8),
    to_signed(-11, 8),
    to_signed(-36, 8),
    to_signed(-59, 8),
    to_signed(-72, 8),
    to_signed(-74, 8),
    to_signed(-64, 8),
    to_signed(-45, 8),
    to_signed(-20, 8),
    to_signed(4, 8),
    to_signed(19, 8),
    to_signed(25, 8),
    to_signed(24, 8),
    to_signed(18, 8),
    to_signed(8, 8),
    to_signed(-4, 8),
    to_signed(-11, 8),
    to_signed(-10, 8),
    to_signed(1, 8),
    to_signed(18, 8),
    to_signed(37, 8),
    to_signed(51, 8),
    to_signed(55, 8),
    to_signed(46, 8),
    to_signed(25, 8),
    to_signed(-1, 8),
    to_signed(-25, 8),
    to_signed(-42, 8),
    to_signed(-51, 8),
    to_signed(-57, 8),
    to_signed(-58, 8),
    to_signed(-56, 8),
    to_signed(-50, 8),
    to_signed(-44, 8),
    to_signed(-42, 8),
    to_signed(-43, 8),
    to_signed(-47, 8),
    to_signed(-53, 8),
    to_signed(-61, 8),
    to_signed(-65, 8),
    to_signed(-62, 8),
    to_signed(-53, 8),
    to_signed(-43, 8),
    to_signed(-34, 8),
    to_signed(-24, 8),
    to_signed(-12, 8),
    to_signed(0, 8),
    to_signed(13, 8),
    to_signed(23, 8),
    to_signed(30, 8),
    to_signed(34, 8),
    to_signed(37, 8),
    to_signed(41, 8),
    to_signed(46, 8),
    to_signed(51, 8),
    to_signed(54, 8),
    to_signed(54, 8),
    to_signed(53, 8),
    to_signed(52, 8),
    to_signed(48, 8),
    to_signed(42, 8),
    to_signed(33, 8),
    to_signed(23, 8),
    to_signed(16, 8),
    to_signed(13, 8),
    to_signed(14, 8),
    to_signed(18, 8),
    to_signed(24, 8),
    to_signed(31, 8),
    to_signed(36, 8),
    to_signed(37, 8),
    to_signed(33, 8),
    to_signed(21, 8),
    to_signed(0, 8),
    to_signed(-29, 8),
    to_signed(-60, 8),
    to_signed(-82, 8),
    to_signed(-89, 8),
    to_signed(-82, 8),
    to_signed(-61, 8),
    to_signed(-34, 8),
    to_signed(-7, 8),
    to_signed(15, 8),
    to_signed(27, 8),
    to_signed(26, 8),
    to_signed(14, 8),
    to_signed(-6, 8),
    to_signed(-27, 8),
    to_signed(-39, 8),
    to_signed(-40, 8),
    to_signed(-28, 8),
    to_signed(-5, 8),
    to_signed(21, 8),
    to_signed(43, 8),
    to_signed(54, 8),
    to_signed(52, 8),
    to_signed(36, 8),
    to_signed(13, 8),
    to_signed(-13, 8),
    to_signed(-37, 8),
    to_signed(-56, 8),
    to_signed(-66, 8),
    to_signed(-65, 8),
    to_signed(-57, 8),
    to_signed(-45, 8),
    to_signed(-36, 8),
    to_signed(-32, 8),
    to_signed(-30, 8),
    to_signed(-32, 8),
    to_signed(-38, 8),
    to_signed(-48, 8),
    to_signed(-56, 8),
    to_signed(-59, 8),
    to_signed(-59, 8),
    to_signed(-55, 8),
    to_signed(-47, 8),
    to_signed(-34, 8),
    to_signed(-19, 8),
    to_signed(-8, 8),
    to_signed(0, 8),
    to_signed(8, 8),
    to_signed(18, 8),
    to_signed(26, 8),
    to_signed(32, 8),
    to_signed(38, 8),
    to_signed(47, 8),
    to_signed(56, 8),
    to_signed(64, 8),
    to_signed(69, 8),
    to_signed(74, 8),
    to_signed(77, 8),
    to_signed(76, 8),
    to_signed(70, 8),
    to_signed(61, 8),
    to_signed(52, 8),
    to_signed(46, 8),
    to_signed(45, 8),
    to_signed(46, 8),
    to_signed(51, 8),
    to_signed(57, 8),
    to_signed(62, 8),
    to_signed(65, 8),
    to_signed(65, 8),
    to_signed(63, 8),
    to_signed(54, 8),
    to_signed(33, 8),
    to_signed(1, 8),
    to_signed(-36, 8),
    to_signed(-69, 8),
    to_signed(-87, 8),
    to_signed(-86, 8),
    to_signed(-67, 8),
    to_signed(-36, 8),
    to_signed(-3, 8),
    to_signed(26, 8),
    to_signed(45, 8),
    to_signed(49, 8),
    to_signed(39, 8),
    to_signed(19, 8),
    to_signed(-6, 8),
    to_signed(-26, 8),
    to_signed(-34, 8),
    to_signed(-28, 8),
    to_signed(-8, 8),
    to_signed(17, 8),
    to_signed(41, 8),
    to_signed(58, 8),
    to_signed(64, 8),
    to_signed(56, 8),
    to_signed(36, 8),
    to_signed(8, 8),
    to_signed(-20, 8),
    to_signed(-44, 8),
    to_signed(-58, 8),
    to_signed(-65, 8),
    to_signed(-64, 8),
    to_signed(-59, 8),
    to_signed(-56, 8),
    to_signed(-53, 8),
    to_signed(-50, 8),
    to_signed(-48, 8),
    to_signed(-48, 8),
    to_signed(-52, 8),
    to_signed(-58, 8),
    to_signed(-61, 8),
    to_signed(-60, 8),
    to_signed(-56, 8),
    to_signed(-50, 8),
    to_signed(-42, 8),
    to_signed(-35, 8),
    to_signed(-27, 8),
    to_signed(-15, 8),
    to_signed(0, 8),
    to_signed(15, 8),
    to_signed(27, 8),
    to_signed(37, 8),
    to_signed(44, 8),
    to_signed(47, 8),
    to_signed(48, 8),
    to_signed(48, 8),
    to_signed(50, 8),
    to_signed(52, 8),
    to_signed(51, 8),
    to_signed(48, 8),
    to_signed(43, 8),
    to_signed(38, 8),
    to_signed(29, 8),
    to_signed(20, 8),
    to_signed(13, 8),
    to_signed(12, 8),
    to_signed(16, 8),
    to_signed(21, 8),
    to_signed(23, 8),
    to_signed(26, 8),
    to_signed(29, 8),
    to_signed(30, 8),
    to_signed(23, 8),
    to_signed(3, 8),
    to_signed(-25, 8),
    to_signed(-55, 8),
    to_signed(-80, 8),
    to_signed(-95, 8),
    to_signed(-92, 8),
    to_signed(-71, 8),
    to_signed(-40, 8),
    to_signed(-9, 8),
    to_signed(19, 8),
    to_signed(39, 8),
    to_signed(47, 8),
    to_signed(41, 8),
    to_signed(24, 8),
    to_signed(2, 8),
    to_signed(-17, 8),
    to_signed(-25, 8),
    to_signed(-20, 8),
    to_signed(-5, 8),
    to_signed(13, 8),
    to_signed(30, 8),
    to_signed(42, 8),
    to_signed(43, 8),
    to_signed(32, 8),
    to_signed(10, 8),
    to_signed(-15, 8),
    to_signed(-38, 8),
    to_signed(-57, 8),
    to_signed(-71, 8),
    to_signed(-79, 8),
    to_signed(-80, 8),
    to_signed(-76, 8),
    to_signed(-70, 8),
    to_signed(-63, 8),
    to_signed(-56, 8),
    to_signed(-52, 8),
    to_signed(-52, 8),
    to_signed(-54, 8),
    to_signed(-54, 8),
    to_signed(-49, 8),
    to_signed(-40, 8),
    to_signed(-33, 8),
    to_signed(-29, 8),
    to_signed(-26, 8),
    to_signed(-21, 8),
    to_signed(-10, 8),
    to_signed(4, 8),
    to_signed(19, 8),
    to_signed(33, 8),
    to_signed(44, 8),
    to_signed(54, 8),
    to_signed(62, 8),
    to_signed(66, 8),
    to_signed(63, 8),
    to_signed(58, 8),
    to_signed(50, 8),
    to_signed(41, 8),
    to_signed(33, 8),
    to_signed(29, 8),
    to_signed(26, 8),
    to_signed(20, 8),
    to_signed(10, 8),
    to_signed(0, 8),
    to_signed(-6, 8),
    to_signed(-6, 8),
    to_signed(-1, 8),
    to_signed(7, 8),
    to_signed(14, 8),
    to_signed(22, 8),
    to_signed(30, 8),
    to_signed(35, 8),
    to_signed(32, 8),
    to_signed(17, 8),
    to_signed(-8, 8),
    to_signed(-38, 8),
    to_signed(-64, 8),
    to_signed(-78, 8),
    to_signed(-78, 8),
    to_signed(-64, 8),
    to_signed(-40, 8),
    to_signed(-12, 8),
    to_signed(16, 8),
    to_signed(40, 8),
    to_signed(53, 8),
    to_signed(52, 8),
    to_signed(39, 8),
    to_signed(20, 8),
    to_signed(-1, 8),
    to_signed(-17, 8),
    to_signed(-21, 8),
    to_signed(-14, 8),
    to_signed(-1, 8),
    to_signed(11, 8),
    to_signed(18, 8),
    to_signed(23, 8),
    to_signed(21, 8),
    to_signed(11, 8),
    to_signed(-7, 8),
    to_signed(-29, 8),
    to_signed(-49, 8),
    to_signed(-64, 8),
    to_signed(-73, 8),
    to_signed(-76, 8),
    to_signed(-73, 8),
    to_signed(-64, 8),
    to_signed(-53, 8),
    to_signed(-44, 8),
    to_signed(-40, 8),
    to_signed(-40, 8),
    to_signed(-39, 8),
    to_signed(-32, 8),
    to_signed(-22, 8),
    to_signed(-12, 8),
    to_signed(-5, 8),
    to_signed(0, 8),
    to_signed(2, 8),
    to_signed(4, 8),
    to_signed(8, 8),
    to_signed(18, 8),
    to_signed(29, 8),
    to_signed(38, 8),
    to_signed(45, 8),
    to_signed(53, 8),
    to_signed(62, 8),
    to_signed(69, 8),
    to_signed(70, 8),
    to_signed(67, 8),
    to_signed(59, 8),
    to_signed(51, 8),
    to_signed(44, 8),
    to_signed(41, 8),
    to_signed(40, 8),
    to_signed(38, 8),
    to_signed(36, 8),
    to_signed(31, 8),
    to_signed(29, 8),
    to_signed(31, 8),
    to_signed(37, 8),
    to_signed(45, 8),
    to_signed(50, 8),
    to_signed(54, 8),
    to_signed(59, 8),
    to_signed(61, 8),
    to_signed(56, 8),
    to_signed(38, 8),
    to_signed(10, 8),
    to_signed(-24, 8),
    to_signed(-56, 8),
    to_signed(-78, 8),
    to_signed(-85, 8),
    to_signed(-75, 8),
    to_signed(-50, 8),
    to_signed(-20, 8),
    to_signed(7, 8),
    to_signed(26, 8),
    to_signed(31, 8),
    to_signed(25, 8),
    to_signed(10, 8),
    to_signed(-9, 8),
    to_signed(-25, 8),
    to_signed(-34, 8),
    to_signed(-32, 8),
    to_signed(-22, 8),
    to_signed(-9, 8),
    to_signed(4, 8),
    to_signed(14, 8),
    to_signed(21, 8),
    to_signed(21, 8),
    to_signed(12, 8),
    to_signed(-4, 8),
    to_signed(-21, 8),
    to_signed(-34, 8),
    to_signed(-43, 8),
    to_signed(-49, 8),
    to_signed(-51, 8),
    to_signed(-48, 8),
    to_signed(-43, 8),
    to_signed(-39, 8),
    to_signed(-36, 8),
    to_signed(-34, 8),
    to_signed(-34, 8),
    to_signed(-33, 8),
    to_signed(-27, 8),
    to_signed(-19, 8),
    to_signed(-14, 8),
    to_signed(-14, 8),
    to_signed(-18, 8),
    to_signed(-25, 8),
    to_signed(-29, 8),
    to_signed(-25, 8),
    to_signed(-14, 8),
    to_signed(0, 8),
    to_signed(11, 8),
    to_signed(23, 8),
    to_signed(36, 8),
    to_signed(48, 8),
    to_signed(56, 8),
    to_signed(59, 8),
    to_signed(56, 8),
    to_signed(48, 8),
    to_signed(40, 8),
    to_signed(35, 8),
    to_signed(35, 8),
    to_signed(37, 8),
    to_signed(38, 8),
    to_signed(38, 8),
    to_signed(38, 8),
    to_signed(40, 8),
    to_signed(44, 8),
    to_signed(48, 8),
    to_signed(52, 8),
    to_signed(52, 8),
    to_signed(50, 8),
    to_signed(46, 8),
    to_signed(35, 8),
    to_signed(16, 8),
    to_signed(-12, 8),
    to_signed(-42, 8),
    to_signed(-70, 8),
    to_signed(-89, 8),
    to_signed(-92, 8),
    to_signed(-78, 8),
    to_signed(-51, 8),
    to_signed(-23, 8),
    to_signed(1, 8),
    to_signed(16, 8),
    to_signed(21, 8),
    to_signed(15, 8),
    to_signed(1, 8),
    to_signed(-16, 8),
    to_signed(-26, 8),
    to_signed(-27, 8),
    to_signed(-19, 8),
    to_signed(-4, 8),
    to_signed(16, 8),
    to_signed(36, 8),
    to_signed(52, 8),
    to_signed(59, 8),
    to_signed(57, 8),
    to_signed(45, 8),
    to_signed(28, 8),
    to_signed(10, 8),
    to_signed(-5, 8),
    to_signed(-17, 8),
    to_signed(-26, 8),
    to_signed(-33, 8),
    to_signed(-38, 8),
    to_signed(-42, 8),
    to_signed(-43, 8),
    to_signed(-42, 8),
    to_signed(-38, 8),
    to_signed(-35, 8),
    to_signed(-36, 8),
    to_signed(-38, 8),
    to_signed(-41, 8),
    to_signed(-43, 8),
    to_signed(-46, 8),
    to_signed(-49, 8),
    to_signed(-48, 8),
    to_signed(-43, 8),
    to_signed(-32, 8),
    to_signed(-13, 8),
    to_signed(10, 8),
    to_signed(31, 8),
    to_signed(49, 8),
    to_signed(62, 8),
    to_signed(72, 8),
    to_signed(76, 8),
    to_signed(75, 8),
    to_signed(69, 8),
    to_signed(60, 8),
    to_signed(51, 8),
    to_signed(45, 8),
    to_signed(42, 8),
    to_signed(41, 8),
    to_signed(42, 8),
    to_signed(44, 8),
    to_signed(49, 8),
    to_signed(54, 8),
    to_signed(57, 8),
    to_signed(55, 8),
    to_signed(48, 8),
    to_signed(39, 8),
    to_signed(26, 8),
    to_signed(9, 8),
    to_signed(-10, 8),
    to_signed(-31, 8),
    to_signed(-51, 8),
    to_signed(-70, 8),
    to_signed(-83, 8),
    to_signed(-84, 8),
    to_signed(-71, 8),
    to_signed(-47, 8),
    to_signed(-21, 8),
    to_signed(0, 8),
    to_signed(12, 8),
    to_signed(14, 8),
    to_signed(9, 8),
    to_signed(-1, 8),
    to_signed(-12, 8),
    to_signed(-19, 8),
    to_signed(-16, 8),
    to_signed(-4, 8),
    to_signed(14, 8),
    to_signed(31, 8),
    to_signed(46, 8),
    to_signed(56, 8),
    to_signed(60, 8),
    to_signed(54, 8),
    to_signed(42, 8),
    to_signed(26, 8),
    to_signed(6, 8),
    to_signed(-16, 8),
    to_signed(-34, 8),
    to_signed(-47, 8),
    to_signed(-53, 8),
    to_signed(-54, 8),
    to_signed(-53, 8),
    to_signed(-51, 8),
    to_signed(-50, 8),
    to_signed(-49, 8),
    to_signed(-50, 8),
    to_signed(-52, 8),
    to_signed(-55, 8),
    to_signed(-57, 8),
    to_signed(-59, 8),
    to_signed(-61, 8),
    to_signed(-61, 8),
    to_signed(-58, 8),
    to_signed(-49, 8),
    to_signed(-33, 8),
    to_signed(-12, 8),
    to_signed(12, 8),
    to_signed(38, 8),
    to_signed(60, 8),
    to_signed(74, 8),
    to_signed(80, 8),
    to_signed(81, 8),
    to_signed(79, 8),
    to_signed(73, 8),
    to_signed(63, 8),
    to_signed(52, 8),
    to_signed(43, 8),
    to_signed(36, 8),
    to_signed(30, 8),
    to_signed(26, 8),
    to_signed(23, 8),
    to_signed(25, 8),
    to_signed(33, 8),
    to_signed(43, 8),
    to_signed(50, 8),
    to_signed(50, 8),
    to_signed(41, 8),
    to_signed(25, 8),
    to_signed(5, 8),
    to_signed(-16, 8),
    to_signed(-37, 8),
    to_signed(-56, 8),
    to_signed(-72, 8),
    to_signed(-83, 8),
    to_signed(-84, 8),
    to_signed(-73, 8),
    to_signed(-51, 8),
    to_signed(-23, 8),
    to_signed(3, 8),
    to_signed(20, 8),
    to_signed(26, 8),
    to_signed(23, 8),
    to_signed(12, 8),
    to_signed(-1, 8),
    to_signed(-12, 8),
    to_signed(-17, 8),
    to_signed(-12, 8),
    to_signed(1, 8),
    to_signed(19, 8),
    to_signed(39, 8),
    to_signed(56, 8),
    to_signed(66, 8),
    to_signed(64, 8),
    to_signed(51, 8),
    to_signed(29, 8),
    to_signed(3, 8),
    to_signed(-21, 8),
    to_signed(-42, 8),
    to_signed(-59, 8),
    to_signed(-68, 8),
    to_signed(-69, 8),
    to_signed(-63, 8),
    to_signed(-55, 8),
    to_signed(-46, 8),
    to_signed(-40, 8),
    to_signed(-38, 8),
    to_signed(-42, 8),
    to_signed(-49, 8),
    to_signed(-54, 8),
    to_signed(-54, 8),
    to_signed(-50, 8),
    to_signed(-43, 8),
    to_signed(-35, 8),
    to_signed(-25, 8),
    to_signed(-12, 8),
    to_signed(5, 8),
    to_signed(25, 8),
    to_signed(45, 8),
    to_signed(62, 8),
    to_signed(74, 8),
    to_signed(78, 8),
    to_signed(76, 8),
    to_signed(70, 8),
    to_signed(63, 8),
    to_signed(54, 8),
    to_signed(46, 8),
    to_signed(38, 8),
    to_signed(33, 8),
    to_signed(29, 8),
    to_signed(23, 8),
    to_signed(16, 8),
    to_signed(10, 8),
    to_signed(7, 8),
    to_signed(9, 8),
    to_signed(14, 8),
    to_signed(18, 8),
    to_signed(18, 8),
    to_signed(15, 8),
    to_signed(9, 8),
    to_signed(3, 8),
    to_signed(-2, 8),
    to_signed(-10, 8),
    to_signed(-22, 8),
    to_signed(-41, 8),
    to_signed(-60, 8),
    to_signed(-72, 8),
    to_signed(-72, 8),
    to_signed(-58, 8),
    to_signed(-35, 8),
    to_signed(-7, 8),
    to_signed(17, 8),
    to_signed(32, 8),
    to_signed(36, 8),
    to_signed(29, 8),
    to_signed(14, 8),
    to_signed(-4, 8),
    to_signed(-19, 8),
    to_signed(-25, 8),
    to_signed(-22, 8),
    to_signed(-12, 8),
    to_signed(3, 8),
    to_signed(18, 8),
    to_signed(30, 8),
    to_signed(36, 8),
    to_signed(33, 8),
    to_signed(20, 8),
    to_signed(-2, 8),
    to_signed(-28, 8),
    to_signed(-50, 8),
    to_signed(-67, 8),
    to_signed(-75, 8),
    to_signed(-75, 8),
    to_signed(-68, 8),
    to_signed(-58, 8),
    to_signed(-50, 8),
    to_signed(-46, 8),
    to_signed(-46, 8),
    to_signed(-49, 8),
    to_signed(-53, 8),
    to_signed(-54, 8),
    to_signed(-52, 8),
    to_signed(-45, 8),
    to_signed(-36, 8),
    to_signed(-28, 8),
    to_signed(-21, 8),
    to_signed(-15, 8),
    to_signed(-7, 8),
    to_signed(3, 8),
    to_signed(17, 8),
    to_signed(31, 8),
    to_signed(44, 8),
    to_signed(54, 8),
    to_signed(60, 8),
    to_signed(63, 8),
    to_signed(64, 8),
    to_signed(60, 8),
    to_signed(54, 8),
    to_signed(48, 8),
    to_signed(41, 8),
    to_signed(33, 8),
    to_signed(25, 8),
    to_signed(18, 8),
    to_signed(12, 8),
    to_signed(9, 8),
    to_signed(9, 8),
    to_signed(13, 8),
    to_signed(22, 8),
    to_signed(29, 8),
    to_signed(31, 8),
    to_signed(29, 8),
    to_signed(25, 8),
    to_signed(22, 8),
    to_signed(18, 8),
    to_signed(7, 8),
    to_signed(-13, 8),
    to_signed(-38, 8),
    to_signed(-60, 8),
    to_signed(-74, 8),
    to_signed(-75, 8),
    to_signed(-64, 8),
    to_signed(-42, 8),
    to_signed(-15, 8),
    to_signed(10, 8),
    to_signed(29, 8),
    to_signed(38, 8),
    to_signed(35, 8),
    to_signed(21, 8),
    to_signed(0, 8),
    to_signed(-20, 8),
    to_signed(-31, 8),
    to_signed(-29, 8),
    to_signed(-17, 8),
    to_signed(-2, 8),
    to_signed(12, 8),
    to_signed(25, 8),
    to_signed(34, 8),
    to_signed(35, 8),
    to_signed(27, 8),
    to_signed(11, 8),
    to_signed(-11, 8),
    to_signed(-30, 8),
    to_signed(-44, 8),
    to_signed(-50, 8),
    to_signed(-50, 8),
    to_signed(-47, 8),
    to_signed(-43, 8),
    to_signed(-42, 8),
    to_signed(-43, 8),
    to_signed(-47, 8),
    to_signed(-48, 8),
    to_signed(-46, 8),
    to_signed(-39, 8),
    to_signed(-31, 8),
    to_signed(-25, 8),
    to_signed(-21, 8),
    to_signed(-20, 8),
    to_signed(-19, 8),
    to_signed(-16, 8),
    to_signed(-10, 8),
    to_signed(-1, 8),
    to_signed(10, 8),
    to_signed(23, 8),
    to_signed(36, 8),
    to_signed(48, 8),
    to_signed(58, 8),
    to_signed(63, 8),
    to_signed(63, 8),
    to_signed(61, 8),
    to_signed(58, 8),
    to_signed(53, 8),
    to_signed(48, 8),
    to_signed(42, 8),
    to_signed(37, 8),
    to_signed(34, 8),
    to_signed(34, 8),
    to_signed(37, 8),
    to_signed(40, 8),
    to_signed(45, 8),
    to_signed(49, 8),
    to_signed(48, 8),
    to_signed(44, 8),
    to_signed(41, 8),
    to_signed(40, 8),
    to_signed(37, 8),
    to_signed(27, 8),
    to_signed(7, 8),
    to_signed(-21, 8),
    to_signed(-50, 8),
    to_signed(-74, 8),
    to_signed(-85, 8),
    to_signed(-82, 8),
    to_signed(-67, 8),
    to_signed(-43, 8),
    to_signed(-16, 8),
    to_signed(10, 8),
    to_signed(27, 8),
    to_signed(32, 8),
    to_signed(24, 8),
    to_signed(8, 8),
    to_signed(-12, 8),
    to_signed(-26, 8),
    to_signed(-30, 8),
    to_signed(-22, 8),
    to_signed(-7, 8),
    to_signed(10, 8),
    to_signed(26, 8),
    to_signed(38, 8),
    to_signed(45, 8),
    to_signed(43, 8),
    to_signed(29, 8),
    to_signed(6, 8),
    to_signed(-18, 8),
    to_signed(-36, 8),
    to_signed(-44, 8),
    to_signed(-46, 8),
    to_signed(-45, 8),
    to_signed(-45, 8),
    to_signed(-46, 8),
    to_signed(-49, 8),
    to_signed(-54, 8),
    to_signed(-59, 8),
    to_signed(-60, 8),
    to_signed(-54, 8),
    to_signed(-43, 8),
    to_signed(-31, 8),
    to_signed(-24, 8),
    to_signed(-24, 8),
    to_signed(-28, 8),
    to_signed(-33, 8),
    to_signed(-34, 8),
    to_signed(-28, 8),
    to_signed(-16, 8),
    to_signed(3, 8),
    to_signed(24, 8),
    to_signed(46, 8),
    to_signed(64, 8),
    to_signed(75, 8),
    to_signed(79, 8),
    to_signed(74, 8),
    to_signed(64, 8),
    to_signed(52, 8),
    to_signed(43, 8),
    to_signed(37, 8),
    to_signed(33, 8),
    to_signed(30, 8),
    to_signed(29, 8),
    to_signed(30, 8),
    to_signed(34, 8),
    to_signed(38, 8),
    to_signed(41, 8),
    to_signed(38, 8),
    to_signed(32, 8),
    to_signed(25, 8),
    to_signed(20, 8),
    to_signed(16, 8),
    to_signed(8, 8),
    to_signed(-7, 8),
    to_signed(-27, 8),
    to_signed(-51, 8),
    to_signed(-71, 8),
    to_signed(-81, 8),
    to_signed(-78, 8),
    to_signed(-64, 8),
    to_signed(-41, 8),
    to_signed(-16, 8),
    to_signed(7, 8),
    to_signed(23, 8),
    to_signed(28, 8),
    to_signed(20, 8),
    to_signed(4, 8),
    to_signed(-13, 8),
    to_signed(-24, 8),
    to_signed(-24, 8),
    to_signed(-14, 8),
    to_signed(3, 8),
    to_signed(22, 8),
    to_signed(37, 8),
    to_signed(46, 8),
    to_signed(49, 8),
    to_signed(44, 8),
    to_signed(30, 8),
    to_signed(8, 8),
    to_signed(-17, 8),
    to_signed(-39, 8),
    to_signed(-53, 8),
    to_signed(-59, 8),
    to_signed(-59, 8),
    to_signed(-57, 8),
    to_signed(-56, 8),
    to_signed(-56, 8),
    to_signed(-59, 8),
    to_signed(-62, 8),
    to_signed(-64, 8),
    to_signed(-63, 8),
    to_signed(-57, 8),
    to_signed(-48, 8),
    to_signed(-40, 8),
    to_signed(-35, 8),
    to_signed(-33, 8),
    to_signed(-30, 8),
    to_signed(-22, 8),
    to_signed(-9, 8),
    to_signed(8, 8),
    to_signed(27, 8),
    to_signed(45, 8),
    to_signed(62, 8),
    to_signed(75, 8),
    to_signed(84, 8),
    to_signed(84, 8),
    to_signed(77, 8),
    to_signed(64, 8),
    to_signed(49, 8),
    to_signed(40, 8),
    to_signed(36, 8),
    to_signed(35, 8),
    to_signed(35, 8),
    to_signed(34, 8),
    to_signed(33, 8),
    to_signed(33, 8),
    to_signed(34, 8),
    to_signed(33, 8),
    to_signed(31, 8),
    to_signed(28, 8),
    to_signed(25, 8),
    to_signed(22, 8),
    to_signed(19, 8),
    to_signed(10, 8),
    to_signed(-6, 8),
    to_signed(-28, 8),
    to_signed(-51, 8),
    to_signed(-71, 8),
    to_signed(-81, 8),
    to_signed(-80, 8),
    to_signed(-66, 8),
    to_signed(-42, 8),
    to_signed(-12, 8),
    to_signed(17, 8),
    to_signed(37, 8),
    to_signed(44, 8),
    to_signed(36, 8),
    to_signed(17, 8),
    to_signed(-4, 8),
    to_signed(-20, 8),
    to_signed(-26, 8),
    to_signed(-21, 8),
    to_signed(-8, 8),
    to_signed(10, 8),
    to_signed(27, 8),
    to_signed(39, 8),
    to_signed(45, 8),
    to_signed(42, 8),
    to_signed(28, 8),
    to_signed(7, 8),
    to_signed(-19, 8),
    to_signed(-43, 8),
    to_signed(-61, 8),
    to_signed(-70, 8),
    to_signed(-71, 8),
    to_signed(-66, 8),
    to_signed(-60, 8),
    to_signed(-56, 8),
    to_signed(-56, 8),
    to_signed(-58, 8),
    to_signed(-60, 8),
    to_signed(-58, 8),
    to_signed(-51, 8),
    to_signed(-41, 8),
    to_signed(-31, 8),
    to_signed(-25, 8),
    to_signed(-23, 8),
    to_signed(-22, 8),
    to_signed(-17, 8),
    to_signed(-7, 8),
    to_signed(6, 8),
    to_signed(22, 8),
    to_signed(38, 8),
    to_signed(52, 8),
    to_signed(63, 8),
    to_signed(72, 8),
    to_signed(76, 8),
    to_signed(72, 8),
    to_signed(61, 8),
    to_signed(46, 8),
    to_signed(34, 8),
    to_signed(26, 8),
    to_signed(24, 8),
    to_signed(24, 8),
    to_signed(26, 8),
    to_signed(30, 8),
    to_signed(35, 8),
    to_signed(39, 8),
    to_signed(41, 8),
    to_signed(39, 8),
    to_signed(34, 8),
    to_signed(29, 8),
    to_signed(25, 8),
    to_signed(21, 8),
    to_signed(14, 8),
    to_signed(3, 8),
    to_signed(-16, 8),
    to_signed(-37, 8),
    to_signed(-57, 8),
    to_signed(-69, 8),
    to_signed(-71, 8),
    to_signed(-62, 8),
    to_signed(-45, 8),
    to_signed(-21, 8),
    to_signed(6, 8),
    to_signed(28, 8),
    to_signed(39, 8),
    to_signed(36, 8),
    to_signed(19, 8),
    to_signed(-3, 8),
    to_signed(-21, 8),
    to_signed(-32, 8),
    to_signed(-31, 8),
    to_signed(-22, 8),
    to_signed(-5, 8),
    to_signed(15, 8),
    to_signed(33, 8),
    to_signed(42, 8),
    to_signed(42, 8),
    to_signed(32, 8),
    to_signed(15, 8),
    to_signed(-7, 8),
    to_signed(-29, 8),
    to_signed(-45, 8),
    to_signed(-54, 8),
    to_signed(-55, 8),
    to_signed(-52, 8),
    to_signed(-48, 8),
    to_signed(-46, 8),
    to_signed(-48, 8),
    to_signed(-51, 8),
    to_signed(-54, 8),
    to_signed(-53, 8),
    to_signed(-49, 8),
    to_signed(-41, 8),
    to_signed(-33, 8),
    to_signed(-29, 8),
    to_signed(-28, 8),
    to_signed(-28, 8),
    to_signed(-24, 8),
    to_signed(-16, 8),
    to_signed(-4, 8),
    to_signed(10, 8),
    to_signed(24, 8),
    to_signed(37, 8),
    to_signed(50, 8),
    to_signed(62, 8),
    to_signed(69, 8),
    to_signed(70, 8),
    to_signed(64, 8),
    to_signed(54, 8),
    to_signed(43, 8),
    to_signed(35, 8),
    to_signed(31, 8),
    to_signed(29, 8),
    to_signed(29, 8),
    to_signed(32, 8),
    to_signed(35, 8),
    to_signed(39, 8),
    to_signed(42, 8),
    to_signed(43, 8),
    to_signed(41, 8),
    to_signed(38, 8),
    to_signed(34, 8),
    to_signed(29, 8),
    to_signed(21, 8),
    to_signed(6, 8),
    to_signed(-17, 8),
    to_signed(-42, 8),
    to_signed(-64, 8),
    to_signed(-77, 8),
    to_signed(-78, 8),
    to_signed(-66, 8),
    to_signed(-43, 8),
    to_signed(-15, 8),
    to_signed(13, 8),
    to_signed(32, 8),
    to_signed(39, 8),
    to_signed(33, 8),
    to_signed(17, 8),
    to_signed(-3, 8),
    to_signed(-21, 8),
    to_signed(-30, 8),
    to_signed(-28, 8),
    to_signed(-17, 8),
    to_signed(3, 8),
    to_signed(25, 8),
    to_signed(44, 8),
    to_signed(55, 8),
    to_signed(56, 8),
    to_signed(46, 8),
    to_signed(26, 8),
    to_signed(-1, 8),
    to_signed(-27, 8),
    to_signed(-46, 8),
    to_signed(-56, 8),
    to_signed(-56, 8),
    to_signed(-51, 8),
    to_signed(-46, 8),
    to_signed(-44, 8),
    to_signed(-47, 8),
    to_signed(-53, 8),
    to_signed(-57, 8),
    to_signed(-57, 8),
    to_signed(-52, 8),
    to_signed(-45, 8),
    to_signed(-37, 8),
    to_signed(-32, 8),
    to_signed(-30, 8),
    to_signed(-30, 8),
    to_signed(-27, 8),
    to_signed(-19, 8),
    to_signed(-6, 8),
    to_signed(8, 8),
    to_signed(21, 8),
    to_signed(32, 8),
    to_signed(41, 8),
    to_signed(50, 8),
    to_signed(57, 8),
    to_signed(58, 8),
    to_signed(54, 8),
    to_signed(46, 8),
    to_signed(39, 8),
    to_signed(33, 8),
    to_signed(31, 8),
    to_signed(32, 8),
    to_signed(34, 8),
    to_signed(36, 8),
    to_signed(38, 8),
    to_signed(40, 8),
    to_signed(41, 8),
    to_signed(39, 8),
    to_signed(33, 8),
    to_signed(24, 8),
    to_signed(12, 8),
    to_signed(1, 8),
    to_signed(-11, 8),
    to_signed(-25, 8),
    to_signed(-40, 8),
    to_signed(-56, 8),
    to_signed(-67, 8),
    to_signed(-70, 8),
    to_signed(-63, 8),
    to_signed(-47, 8),
    to_signed(-24, 8),
    to_signed(1, 8),
    to_signed(21, 8),
    to_signed(34, 8),
    to_signed(36, 8),
    to_signed(28, 8),
    to_signed(13, 8),
    to_signed(-4, 8),
    to_signed(-16, 8),
    to_signed(-18, 8),
    to_signed(-10, 8),
    to_signed(6, 8),
    to_signed(26, 8),
    to_signed(44, 8),
    to_signed(55, 8),
    to_signed(57, 8),
    to_signed(50, 8),
    to_signed(36, 8),
    to_signed(16, 8),
    to_signed(-9, 8),
    to_signed(-32, 8),
    to_signed(-50, 8),
    to_signed(-59, 8),
    to_signed(-59, 8),
    to_signed(-54, 8),
    to_signed(-47, 8),
    to_signed(-44, 8),
    to_signed(-45, 8),
    to_signed(-49, 8),
    to_signed(-52, 8),
    to_signed(-53, 8),
    to_signed(-50, 8),
    to_signed(-43, 8),
    to_signed(-35, 8),
    to_signed(-28, 8),
    to_signed(-25, 8),
    to_signed(-23, 8),
    to_signed(-19, 8),
    to_signed(-11, 8),
    to_signed(3, 8),
    to_signed(19, 8),
    to_signed(34, 8),
    to_signed(47, 8),
    to_signed(58, 8),
    to_signed(66, 8),
    to_signed(69, 8),
    to_signed(67, 8),
    to_signed(60, 8),
    to_signed(50, 8),
    to_signed(39, 8),
    to_signed(31, 8),
    to_signed(27, 8),
    to_signed(27, 8),
    to_signed(29, 8),
    to_signed(30, 8),
    to_signed(31, 8),
    to_signed(31, 8),
    to_signed(31, 8),
    to_signed(31, 8),
    to_signed(29, 8),
    to_signed(23, 8),
    to_signed(15, 8),
    to_signed(6, 8),
    to_signed(-5, 8),
    to_signed(-19, 8),
    to_signed(-38, 8),
    to_signed(-57, 8),
    to_signed(-70, 8),
    to_signed(-72, 8),
    to_signed(-61, 8),
    to_signed(-40, 8),
    to_signed(-14, 8),
    to_signed(11, 8),
    to_signed(31, 8),
    to_signed(42, 8),
    to_signed(44, 8),
    to_signed(37, 8),
    to_signed(21, 8),
    to_signed(3, 8),
    to_signed(-11, 8),
    to_signed(-17, 8),
    to_signed(-12, 8),
    to_signed(2, 8),
    to_signed(21, 8),
    to_signed(38, 8),
    to_signed(49, 8),
    to_signed(53, 8),
    to_signed(47, 8),
    to_signed(33, 8),
    to_signed(11, 8),
    to_signed(-15, 8),
    to_signed(-38, 8),
    to_signed(-56, 8),
    to_signed(-65, 8),
    to_signed(-67, 8),
    to_signed(-64, 8),
    to_signed(-59, 8),
    to_signed(-55, 8),
    to_signed(-54, 8),
    to_signed(-53, 8),
    to_signed(-53, 8),
    to_signed(-52, 8),
    to_signed(-47, 8),
    to_signed(-42, 8),
    to_signed(-35, 8),
    to_signed(-30, 8),
    to_signed(-26, 8),
    to_signed(-22, 8),
    to_signed(-16, 8),
    to_signed(-6, 8),
    to_signed(8, 8),
    to_signed(24, 8),
    to_signed(42, 8),
    to_signed(57, 8),
    to_signed(69, 8),
    to_signed(75, 8),
    to_signed(75, 8),
    to_signed(70, 8),
    to_signed(59, 8),
    to_signed(45, 8),
    to_signed(30, 8),
    to_signed(19, 8),
    to_signed(14, 8),
    to_signed(14, 8),
    to_signed(17, 8),
    to_signed(20, 8),
    to_signed(22, 8),
    to_signed(22, 8),
    to_signed(21, 8),
    to_signed(19, 8),
    to_signed(16, 8),
    to_signed(12, 8),
    to_signed(9, 8),
    to_signed(9, 8),
    to_signed(9, 8),
    to_signed(6, 8),
    to_signed(-4, 8),
    to_signed(-20, 8),
    to_signed(-39, 8),
    to_signed(-55, 8),
    to_signed(-60, 8),
    to_signed(-53, 8),
    to_signed(-36, 8),
    to_signed(-12, 8),
    to_signed(13, 8),
    to_signed(36, 8),
    to_signed(51, 8),
    to_signed(52, 8),
    to_signed(40, 8),
    to_signed(18, 8),
    to_signed(-6, 8),
    to_signed(-26, 8),
    to_signed(-36, 8),
    to_signed(-35, 8),
    to_signed(-25, 8),
    to_signed(-9, 8),
    to_signed(9, 8),
    to_signed(24, 8),
    to_signed(31, 8),
    to_signed(29, 8),
    to_signed(16, 8),
    to_signed(-5, 8),
    to_signed(-31, 8),
    to_signed(-54, 8),
    to_signed(-70, 8),
    to_signed(-75, 8),
    to_signed(-73, 8),
    to_signed(-68, 8),
    to_signed(-62, 8),
    to_signed(-56, 8),
    to_signed(-51, 8),
    to_signed(-46, 8),
    to_signed(-41, 8),
    to_signed(-35, 8),
    to_signed(-29, 8),
    to_signed(-23, 8),
    to_signed(-17, 8),
    to_signed(-15, 8),
    to_signed(-16, 8),
    to_signed(-18, 8),
    to_signed(-17, 8),
    to_signed(-11, 8),
    to_signed(-2, 8),
    to_signed(11, 8),
    to_signed(24, 8),
    to_signed(38, 8),
    to_signed(50, 8),
    to_signed(59, 8),
    to_signed(64, 8),
    to_signed(65, 8),
    to_signed(59, 8),
    to_signed(50, 8),
    to_signed(41, 8),
    to_signed(37, 8),
    to_signed(36, 8),
    to_signed(35, 8),
    to_signed(35, 8),
    to_signed(34, 8),
    to_signed(34, 8),
    to_signed(34, 8),
    to_signed(34, 8),
    to_signed(32, 8),
    to_signed(30, 8),
    to_signed(28, 8),
    to_signed(26, 8),
    to_signed(23, 8),
    to_signed(15, 8),
    to_signed(0, 8),
    to_signed(-22, 8),
    to_signed(-46, 8),
    to_signed(-66, 8),
    to_signed(-77, 8),
    to_signed(-77, 8),
    to_signed(-65, 8),
    to_signed(-42, 8),
    to_signed(-14, 8),
    to_signed(13, 8),
    to_signed(34, 8),
    to_signed(43, 8),
    to_signed(40, 8),
    to_signed(25, 8),
    to_signed(6, 8),
    to_signed(-9, 8),
    to_signed(-15, 8),
    to_signed(-11, 8),
    to_signed(1, 8),
    to_signed(16, 8),
    to_signed(33, 8),
    to_signed(46, 8),
    to_signed(52, 8),
    to_signed(51, 8),
    to_signed(39, 8),
    to_signed(17, 8),
    to_signed(-9, 8),
    to_signed(-33, 8),
    to_signed(-51, 8),
    to_signed(-62, 8),
    to_signed(-69, 8),
    to_signed(-73, 8),
    to_signed(-74, 8),
    to_signed(-73, 8),
    to_signed(-71, 8),
    to_signed(-67, 8),
    to_signed(-62, 8),
    to_signed(-55, 8),
    to_signed(-44, 8),
    to_signed(-32, 8),
    to_signed(-19, 8),
    to_signed(-11, 8),
    to_signed(-8, 8),
    to_signed(-9, 8),
    to_signed(-10, 8),
    to_signed(-7, 8),
    to_signed(1, 8),
    to_signed(13, 8),
    to_signed(28, 8),
    to_signed(45, 8),
    to_signed(60, 8),
    to_signed(72, 8),
    to_signed(79, 8),
    to_signed(78, 8),
    to_signed(69, 8),
    to_signed(55, 8),
    to_signed(41, 8),
    to_signed(28, 8),
    to_signed(18, 8),
    to_signed(10, 8),
    to_signed(7, 8),
    to_signed(8, 8),
    to_signed(13, 8),
    to_signed(18, 8),
    to_signed(22, 8),
    to_signed(25, 8),
    to_signed(24, 8),
    to_signed(22, 8),
    to_signed(19, 8),
    to_signed(16, 8),
    to_signed(10, 8),
    to_signed(-1, 8),
    to_signed(-17, 8),
    to_signed(-35, 8),
    to_signed(-53, 8),
    to_signed(-64, 8),
    to_signed(-66, 8),
    to_signed(-57, 8),
    to_signed(-37, 8),
    to_signed(-11, 8),
    to_signed(17, 8),
    to_signed(40, 8),
    to_signed(52, 8),
    to_signed(50, 8),
    to_signed(37, 8),
    to_signed(17, 8),
    to_signed(-2, 8),
    to_signed(-16, 8),
    to_signed(-23, 8),
    to_signed(-22, 8),
    to_signed(-14, 8),
    to_signed(0, 8),
    to_signed(14, 8),
    to_signed(25, 8),
    to_signed(29, 8),
    to_signed(22, 8),
    to_signed(5, 8),
    to_signed(-17, 8),
    to_signed(-37, 8),
    to_signed(-51, 8),
    to_signed(-60, 8),
    to_signed(-65, 8),
    to_signed(-68, 8),
    to_signed(-69, 8),
    to_signed(-67, 8),
    to_signed(-65, 8),
    to_signed(-62, 8),
    to_signed(-57, 8),
    to_signed(-48, 8),
    to_signed(-36, 8),
    to_signed(-21, 8),
    to_signed(-8, 8),
    to_signed(-1, 8),
    to_signed(-2, 8),
    to_signed(-7, 8),
    to_signed(-13, 8),
    to_signed(-15, 8),
    to_signed(-11, 8),
    to_signed(0, 8),
    to_signed(16, 8),
    to_signed(37, 8),
    to_signed(59, 8),
    to_signed(77, 8),
    to_signed(87, 8),
    to_signed(86, 8),
    to_signed(75, 8),
    to_signed(59, 8),
    to_signed(42, 8),
    to_signed(29, 8),
    to_signed(21, 8),
    to_signed(19, 8),
    to_signed(21, 8),
    to_signed(25, 8),
    to_signed(29, 8),
    to_signed(33, 8),
    to_signed(36, 8),
    to_signed(37, 8),
    to_signed(37, 8),
    to_signed(35, 8),
    to_signed(33, 8),
    to_signed(30, 8),
    to_signed(24, 8),
    to_signed(11, 8),
    to_signed(-9, 8),
    to_signed(-36, 8),
    to_signed(-62, 8),
    to_signed(-83, 8),
    to_signed(-93, 8),
    to_signed(-89, 8),
    to_signed(-69, 8),
    to_signed(-39, 8),
    to_signed(-7, 8),
    to_signed(19, 8),
    to_signed(32, 8),
    to_signed(31, 8),
    to_signed(19, 8),
    to_signed(2, 8),
    to_signed(-13, 8),
    to_signed(-22, 8),
    to_signed(-23, 8),
    to_signed(-17, 8),
    to_signed(-4, 8),
    to_signed(11, 8),
    to_signed(25, 8),
    to_signed(33, 8),
    to_signed(34, 8),
    to_signed(27, 8),
    to_signed(12, 8),
    to_signed(-6, 8),
    to_signed(-24, 8),
    to_signed(-39, 8),
    to_signed(-50, 8),
    to_signed(-57, 8),
    to_signed(-60, 8),
    to_signed(-61, 8),
    to_signed(-63, 8),
    to_signed(-66, 8),
    to_signed(-68, 8),
    to_signed(-63, 8),
    to_signed(-52, 8),
    to_signed(-37, 8),
    to_signed(-22, 8),
    to_signed(-12, 8),
    to_signed(-7, 8),
    to_signed(-8, 8),
    to_signed(-12, 8),
    to_signed(-16, 8),
    to_signed(-13, 8),
    to_signed(-4, 8),
    to_signed(10, 8),
    to_signed(27, 8),
    to_signed(44, 8),
    to_signed(60, 8),
    to_signed(72, 8),
    to_signed(77, 8),
    to_signed(75, 8),
    to_signed(67, 8),
    to_signed(55, 8),
    to_signed(43, 8),
    to_signed(35, 8),
    to_signed(30, 8),
    to_signed(26, 8),
    to_signed(23, 8),
    to_signed(23, 8),
    to_signed(25, 8),
    to_signed(27, 8),
    to_signed(29, 8),
    to_signed(30, 8),
    to_signed(29, 8),
    to_signed(25, 8),
    to_signed(19, 8),
    to_signed(12, 8),
    to_signed(3, 8),
    to_signed(-10, 8),
    to_signed(-27, 8),
    to_signed(-45, 8),
    to_signed(-59, 8),
    to_signed(-67, 8),
    to_signed(-66, 8),
    to_signed(-55, 8),
    to_signed(-34, 8),
    to_signed(-8, 8),
    to_signed(15, 8),
    to_signed(33, 8),
    to_signed(40, 8),
    to_signed(37, 8),
    to_signed(27, 8),
    to_signed(14, 8),
    to_signed(3, 8),
    to_signed(-4, 8),
    to_signed(-5, 8),
    to_signed(0, 8),
    to_signed(10, 8),
    to_signed(18, 8),
    to_signed(22, 8),
    to_signed(21, 8),
    to_signed(17, 8),
    to_signed(10, 8),
    to_signed(-1, 8),
    to_signed(-16, 8),
    to_signed(-30, 8),
    to_signed(-42, 8),
    to_signed(-49, 8),
    to_signed(-52, 8),
    to_signed(-53, 8),
    to_signed(-55, 8),
    to_signed(-59, 8),
    to_signed(-63, 8),
    to_signed(-63, 8),
    to_signed(-57, 8),
    to_signed(-44, 8),
    to_signed(-30, 8),
    to_signed(-16, 8),
    to_signed(-6, 8),
    to_signed(-1, 8),
    to_signed(-1, 8),
    to_signed(-6, 8),
    to_signed(-9, 8),
    to_signed(-9, 8),
    to_signed(-4, 8),
    to_signed(5, 8),
    to_signed(18, 8),
    to_signed(33, 8),
    to_signed(47, 8),
    to_signed(57, 8),
    to_signed(59, 8),
    to_signed(54, 8),
    to_signed(44, 8),
    to_signed(31, 8),
    to_signed(21, 8),
    to_signed(16, 8),
    to_signed(16, 8),
    to_signed(19, 8),
    to_signed(24, 8),
    to_signed(30, 8),
    to_signed(34, 8),
    to_signed(36, 8),
    to_signed(36, 8),
    to_signed(35, 8),
    to_signed(33, 8),
    to_signed(28, 8),
    to_signed(21, 8),
    to_signed(11, 8),
    to_signed(-4, 8),
    to_signed(-23, 8),
    to_signed(-44, 8),
    to_signed(-60, 8),
    to_signed(-69, 8),
    to_signed(-68, 8),
    to_signed(-57, 8),
    to_signed(-37, 8),
    to_signed(-12, 8),
    to_signed(10, 8),
    to_signed(25, 8),
    to_signed(30, 8),
    to_signed(26, 8),
    to_signed(15, 8),
    to_signed(1, 8),
    to_signed(-10, 8),
    to_signed(-14, 8),
    to_signed(-9, 8),
    to_signed(5, 8),
    to_signed(21, 8),
    to_signed(35, 8),
    to_signed(42, 8),
    to_signed(42, 8),
    to_signed(37, 8),
    to_signed(28, 8),
    to_signed(16, 8),
    to_signed(3, 8),
    to_signed(-12, 8),
    to_signed(-26, 8),
    to_signed(-37, 8),
    to_signed(-45, 8),
    to_signed(-50, 8),
    to_signed(-53, 8),
    to_signed(-56, 8),
    to_signed(-57, 8),
    to_signed(-57, 8),
    to_signed(-52, 8),
    to_signed(-40, 8),
    to_signed(-25, 8),
    to_signed(-13, 8),
    to_signed(-7, 8),
    to_signed(-8, 8),
    to_signed(-15, 8),
    to_signed(-24, 8),
    to_signed(-31, 8),
    to_signed(-29, 8),
    to_signed(-18, 8),
    to_signed(0, 8),
    to_signed(22, 8),
    to_signed(42, 8),
    to_signed(59, 8),
    to_signed(69, 8),
    to_signed(71, 8),
    to_signed(67, 8),
    to_signed(59, 8),
    to_signed(48, 8),
    to_signed(35, 8),
    to_signed(23, 8),
    to_signed(13, 8),
    to_signed(9, 8),
    to_signed(9, 8),
    to_signed(14, 8),
    to_signed(21, 8),
    to_signed(27, 8),
    to_signed(29, 8),
    to_signed(29, 8),
    to_signed(26, 8),
    to_signed(21, 8),
    to_signed(12, 8),
    to_signed(0, 8),
    to_signed(-15, 8),
    to_signed(-32, 8),
    to_signed(-49, 8),
    to_signed(-63, 8),
    to_signed(-69, 8),
    to_signed(-63, 8),
    to_signed(-47, 8),
    to_signed(-23, 8),
    to_signed(3, 8),
    to_signed(24, 8),
    to_signed(36, 8),
    to_signed(37, 8),
    to_signed(30, 8),
    to_signed(18, 8),
    to_signed(6, 8),
    to_signed(-4, 8),
    to_signed(-7, 8),
    to_signed(-3, 8),
    to_signed(8, 8),
    to_signed(22, 8),
    to_signed(36, 8),
    to_signed(45, 8),
    to_signed(48, 8),
    to_signed(43, 8),
    to_signed(30, 8),
    to_signed(14, 8),
    to_signed(-2, 8),
    to_signed(-18, 8),
    to_signed(-32, 8),
    to_signed(-43, 8),
    to_signed(-49, 8),
    to_signed(-52, 8),
    to_signed(-51, 8),
    to_signed(-48, 8),
    to_signed(-44, 8),
    to_signed(-41, 8),
    to_signed(-36, 8),
    to_signed(-30, 8),
    to_signed(-22, 8),
    to_signed(-14, 8),
    to_signed(-9, 8),
    to_signed(-9, 8),
    to_signed(-13, 8),
    to_signed(-20, 8),
    to_signed(-25, 8),
    to_signed(-23, 8),
    to_signed(-13, 8),
    to_signed(3, 8),
    to_signed(23, 8),
    to_signed(42, 8),
    to_signed(57, 8),
    to_signed(66, 8),
    to_signed(66, 8),
    to_signed(58, 8),
    to_signed(47, 8),
    to_signed(35, 8),
    to_signed(24, 8),
    to_signed(15, 8),
    to_signed(7, 8),
    to_signed(2, 8),
    to_signed(0, 8),
    to_signed(3, 8),
    to_signed(8, 8),
    to_signed(16, 8),
    to_signed(22, 8),
    to_signed(27, 8),
    to_signed(30, 8),
    to_signed(29, 8),
    to_signed(22, 8),
    to_signed(11, 8),
    to_signed(-4, 8),
    to_signed(-22, 8),
    to_signed(-41, 8),
    to_signed(-60, 8),
    to_signed(-72, 8),
    to_signed(-74, 8),
    to_signed(-64, 8),
    to_signed(-42, 8),
    to_signed(-13, 8),
    to_signed(16, 8),
    to_signed(36, 8),
    to_signed(43, 8),
    to_signed(37, 8),
    to_signed(21, 8),
    to_signed(2, 8),
    to_signed(-15, 8),
    to_signed(-25, 8),
    to_signed(-25, 8),
    to_signed(-16, 8),
    to_signed(-1, 8),
    to_signed(17, 8),
    to_signed(31, 8),
    to_signed(40, 8),
    to_signed(43, 8),
    to_signed(39, 8),
    to_signed(30, 8),
    to_signed(16, 8),
    to_signed(0, 8),
    to_signed(-14, 8),
    to_signed(-26, 8),
    to_signed(-34, 8),
    to_signed(-39, 8),
    to_signed(-41, 8),
    to_signed(-42, 8),
    to_signed(-40, 8),
    to_signed(-39, 8),
    to_signed(-37, 8),
    to_signed(-35, 8),
    to_signed(-31, 8),
    to_signed(-25, 8),
    to_signed(-18, 8),
    to_signed(-14, 8),
    to_signed(-14, 8),
    to_signed(-18, 8),
    to_signed(-24, 8),
    to_signed(-26, 8),
    to_signed(-22, 8),
    to_signed(-11, 8),
    to_signed(4, 8),
    to_signed(19, 8),
    to_signed(33, 8),
    to_signed(44, 8),
    to_signed(51, 8),
    to_signed(53, 8),
    to_signed(51, 8),
    to_signed(44, 8),
    to_signed(35, 8),
    to_signed(25, 8),
    to_signed(15, 8),
    to_signed(8, 8),
    to_signed(3, 8),
    to_signed(3, 8),
    to_signed(7, 8),
    to_signed(14, 8),
    to_signed(22, 8),
    to_signed(30, 8),
    to_signed(35, 8),
    to_signed(37, 8),
    to_signed(34, 8),
    to_signed(27, 8),
    to_signed(17, 8),
    to_signed(3, 8),
    to_signed(-14, 8),
    to_signed(-35, 8),
    to_signed(-57, 8),
    to_signed(-73, 8),
    to_signed(-80, 8),
    to_signed(-73, 8),
    to_signed(-53, 8),
    to_signed(-25, 8),
    to_signed(2, 8),
    to_signed(24, 8),
    to_signed(38, 8),
    to_signed(40, 8),
    to_signed(32, 8),
    to_signed(18, 8),
    to_signed(3, 8),
    to_signed(-7, 8),
    to_signed(-11, 8),
    to_signed(-7, 8),
    to_signed(4, 8),
    to_signed(18, 8),
    to_signed(32, 8),
    to_signed(44, 8),
    to_signed(52, 8),
    to_signed(52, 8),
    to_signed(44, 8),
    to_signed(29, 8),
    to_signed(10, 8),
    to_signed(-7, 8),
    to_signed(-22, 8),
    to_signed(-34, 8),
    to_signed(-42, 8),
    to_signed(-48, 8),
    to_signed(-52, 8),
    to_signed(-55, 8),
    to_signed(-59, 8),
    to_signed(-62, 8),
    to_signed(-62, 8),
    to_signed(-56, 8),
    to_signed(-44, 8),
    to_signed(-29, 8),
    to_signed(-15, 8),
    to_signed(-7, 8),
    to_signed(-6, 8),
    to_signed(-9, 8),
    to_signed(-11, 8),
    to_signed(-10, 8),
    to_signed(-6, 8),
    to_signed(3, 8),
    to_signed(14, 8),
    to_signed(27, 8),
    to_signed(42, 8),
    to_signed(55, 8),
    to_signed(63, 8),
    to_signed(64, 8),
    to_signed(60, 8),
    to_signed(50, 8),
    to_signed(40, 8),
    to_signed(29, 8),
    to_signed(20, 8),
    to_signed(13, 8),
    to_signed(10, 8),
    to_signed(10, 8),
    to_signed(15, 8),
    to_signed(22, 8),
    to_signed(28, 8),
    to_signed(31, 8),
    to_signed(29, 8),
    to_signed(24, 8),
    to_signed(18, 8),
    to_signed(10, 8),
    to_signed(-3, 8),
    to_signed(-19, 8),
    to_signed(-38, 8),
    to_signed(-59, 8),
    to_signed(-76, 8),
    to_signed(-83, 8),
    to_signed(-78, 8),
    to_signed(-62, 8),
    to_signed(-38, 8),
    to_signed(-11, 8),
    to_signed(15, 8),
    to_signed(34, 8),
    to_signed(41, 8),
    to_signed(36, 8),
    to_signed(23, 8),
    to_signed(8, 8),
    to_signed(-5, 8),
    to_signed(-15, 8),
    to_signed(-16, 8),
    to_signed(-10, 8),
    to_signed(2, 8),
    to_signed(15, 8),
    to_signed(27, 8),
    to_signed(38, 8),
    to_signed(44, 8),
    to_signed(40, 8),
    to_signed(29, 8),
    to_signed(12, 8),
    to_signed(-7, 8),
    to_signed(-25, 8),
    to_signed(-39, 8),
    to_signed(-49, 8),
    to_signed(-55, 8),
    to_signed(-59, 8),
    to_signed(-61, 8),
    to_signed(-61, 8),
    to_signed(-59, 8),
    to_signed(-53, 8),
    to_signed(-43, 8),
    to_signed(-31, 8),
    to_signed(-17, 8),
    to_signed(-6, 8),
    to_signed(0, 8),
    to_signed(0, 8),
    to_signed(-5, 8),
    to_signed(-9, 8),
    to_signed(-9, 8),
    to_signed(-6, 8),
    to_signed(2, 8),
    to_signed(13, 8),
    to_signed(26, 8),
    to_signed(41, 8),
    to_signed(56, 8),
    to_signed(65, 8),
    to_signed(66, 8),
    to_signed(60, 8),
    to_signed(49, 8),
    to_signed(35, 8),
    to_signed(22, 8),
    to_signed(13, 8),
    to_signed(8, 8),
    to_signed(7, 8),
    to_signed(11, 8),
    to_signed(18, 8),
    to_signed(26, 8),
    to_signed(30, 8),
    to_signed(31, 8),
    to_signed(30, 8),
    to_signed(28, 8),
    to_signed(23, 8),
    to_signed(11, 8),
    to_signed(-7, 8),
    to_signed(-29, 8),
    to_signed(-51, 8),
    to_signed(-71, 8),
    to_signed(-82, 8),
    to_signed(-81, 8),
    to_signed(-67, 8),
    to_signed(-45, 8),
    to_signed(-17, 8),
    to_signed(11, 8),
    to_signed(34, 8),
    to_signed(45, 8),
    to_signed(44, 8),
    to_signed(33, 8),
    to_signed(17, 8),
    to_signed(1, 8),
    to_signed(-12, 8),
    to_signed(-19, 8),
    to_signed(-16, 8),
    to_signed(-6, 8),
    to_signed(8, 8),
    to_signed(22, 8),
    to_signed(35, 8),
    to_signed(44, 8),
    to_signed(46, 8),
    to_signed(38, 8),
    to_signed(24, 8),
    to_signed(6, 8),
    to_signed(-11, 8),
    to_signed(-25, 8),
    to_signed(-36, 8),
    to_signed(-45, 8),
    to_signed(-51, 8),
    to_signed(-55, 8),
    to_signed(-55, 8),
    to_signed(-51, 8),
    to_signed(-45, 8),
    to_signed(-38, 8),
    to_signed(-29, 8),
    to_signed(-18, 8),
    to_signed(-8, 8),
    to_signed(-3, 8),
    to_signed(-2, 8),
    to_signed(-7, 8),
    to_signed(-14, 8),
    to_signed(-16, 8),
    to_signed(-10, 8),
    to_signed(3, 8),
    to_signed(17, 8),
    to_signed(32, 8),
    to_signed(47, 8),
    to_signed(61, 8),
    to_signed(70, 8),
    to_signed(72, 8),
    to_signed(68, 8),
    to_signed(59, 8),
    to_signed(48, 8),
    to_signed(36, 8),
    to_signed(26, 8),
    to_signed(19, 8),
    to_signed(15, 8),
    to_signed(15, 8),
    to_signed(18, 8),
    to_signed(24, 8),
    to_signed(30, 8),
    to_signed(32, 8),
    to_signed(32, 8),
    to_signed(29, 8),
    to_signed(22, 8),
    to_signed(8, 8),
    to_signed(-14, 8),
    to_signed(-40, 8),
    to_signed(-64, 8),
    to_signed(-83, 8),
    to_signed(-92, 8),
    to_signed(-91, 8),
    to_signed(-77, 8),
    to_signed(-52, 8),
    to_signed(-19, 8),
    to_signed(14, 8),
    to_signed(39, 8),
    to_signed(50, 8),
    to_signed(46, 8),
    to_signed(31, 8),
    to_signed(13, 8),
    to_signed(-4, 8),
    to_signed(-15, 8),
    to_signed(-18, 8),
    to_signed(-13, 8),
    to_signed(-1, 8),
    to_signed(14, 8),
    to_signed(30, 8),
    to_signed(40, 8),
    to_signed(43, 8),
    to_signed(38, 8),
    to_signed(27, 8),
    to_signed(12, 8),
    to_signed(-5, 8),
    to_signed(-20, 8),
    to_signed(-32, 8),
    to_signed(-42, 8),
    to_signed(-50, 8),
    to_signed(-56, 8),
    to_signed(-59, 8),
    to_signed(-59, 8),
    to_signed(-58, 8),
    to_signed(-54, 8),
    to_signed(-47, 8),
    to_signed(-36, 8),
    to_signed(-23, 8),
    to_signed(-12, 8),
    to_signed(-6, 8),
    to_signed(-4, 8),
    to_signed(-7, 8),
    to_signed(-12, 8),
    to_signed(-14, 8),
    to_signed(-8, 8),
    to_signed(5, 8),
    to_signed(22, 8),
    to_signed(37, 8),
    to_signed(49, 8),
    to_signed(58, 8),
    to_signed(62, 8),
    to_signed(58, 8),
    to_signed(48, 8),
    to_signed(35, 8),
    to_signed(19, 8),
    to_signed(3, 8),
    to_signed(-9, 8),
    to_signed(-16, 8),
    to_signed(-17, 8),
    to_signed(-14, 8),
    to_signed(-7, 8),
    to_signed(0, 8),
    to_signed(7, 8),
    to_signed(13, 8),
    to_signed(17, 8),
    to_signed(19, 8),
    to_signed(16, 8),
    to_signed(7, 8),
    to_signed(-7, 8),
    to_signed(-28, 8),
    to_signed(-50, 8),
    to_signed(-70, 8),
    to_signed(-80, 8),
    to_signed(-79, 8),
    to_signed(-66, 8),
    to_signed(-42, 8),
    to_signed(-9, 8),
    to_signed(23, 8),
    to_signed(47, 8),
    to_signed(57, 8),
    to_signed(50, 8),
    to_signed(32, 8),
    to_signed(9, 8),
    to_signed(-11, 8),
    to_signed(-23, 8),
    to_signed(-27, 8),
    to_signed(-22, 8),
    to_signed(-10, 8),
    to_signed(7, 8),
    to_signed(24, 8),
    to_signed(35, 8),
    to_signed(37, 8),
    to_signed(31, 8),
    to_signed(20, 8),
    to_signed(9, 8),
    to_signed(-3, 8),
    to_signed(-15, 8),
    to_signed(-24, 8),
    to_signed(-31, 8),
    to_signed(-38, 8),
    to_signed(-42, 8),
    to_signed(-43, 8),
    to_signed(-42, 8),
    to_signed(-41, 8),
    to_signed(-39, 8),
    to_signed(-34, 8),
    to_signed(-27, 8),
    to_signed(-18, 8),
    to_signed(-10, 8),
    to_signed(-5, 8),
    to_signed(-2, 8),
    to_signed(-3, 8),
    to_signed(-6, 8),
    to_signed(-10, 8),
    to_signed(-9, 8),
    to_signed(-1, 8),
    to_signed(13, 8),
    to_signed(28, 8),
    to_signed(43, 8),
    to_signed(53, 8),
    to_signed(59, 8),
    to_signed(59, 8),
    to_signed(55, 8),
    to_signed(48, 8),
    to_signed(39, 8),
    to_signed(30, 8),
    to_signed(21, 8),
    to_signed(13, 8),
    to_signed(7, 8),
    to_signed(2, 8),
    to_signed(2, 8),
    to_signed(7, 8),
    to_signed(14, 8),
    to_signed(23, 8),
    to_signed(30, 8),
    to_signed(35, 8),
    to_signed(33, 8),
    to_signed(23, 8),
    to_signed(6, 8),
    to_signed(-17, 8),
    to_signed(-44, 8),
    to_signed(-69, 8),
    to_signed(-84, 8),
    to_signed(-87, 8),
    to_signed(-75, 8),
    to_signed(-52, 8),
    to_signed(-20, 8),
    to_signed(13, 8),
    to_signed(38, 8),
    to_signed(51, 8),
    to_signed(49, 8),
    to_signed(33, 8),
    to_signed(11, 8),
    to_signed(-7, 8),
    to_signed(-17, 8),
    to_signed(-17, 8),
    to_signed(-8, 8),
    to_signed(7, 8),
    to_signed(25, 8),
    to_signed(42, 8),
    to_signed(52, 8),
    to_signed(54, 8),
    to_signed(47, 8),
    to_signed(31, 8),
    to_signed(11, 8),
    to_signed(-8, 8),
    to_signed(-23, 8),
    to_signed(-35, 8),
    to_signed(-43, 8),
    to_signed(-48, 8),
    to_signed(-52, 8),
    to_signed(-55, 8),
    to_signed(-56, 8),
    to_signed(-56, 8),
    to_signed(-56, 8),
    to_signed(-52, 8),
    to_signed(-45, 8),
    to_signed(-35, 8),
    to_signed(-28, 8),
    to_signed(-23, 8),
    to_signed(-18, 8),
    to_signed(-13, 8),
    to_signed(-9, 8),
    to_signed(-5, 8),
    to_signed(1, 8),
    to_signed(11, 8),
    to_signed(23, 8),
    to_signed(34, 8),
    to_signed(44, 8),
    to_signed(52, 8),
    to_signed(55, 8),
    to_signed(55, 8),
    to_signed(51, 8),
    to_signed(46, 8),
    to_signed(39, 8),
    to_signed(30, 8),
    to_signed(21, 8),
    to_signed(13, 8),
    to_signed(5, 8),
    to_signed(-2, 8),
    to_signed(-5, 8),
    to_signed(-2, 8),
    to_signed(5, 8),
    to_signed(13, 8),
    to_signed(20, 8),
    to_signed(26, 8),
    to_signed(26, 8),
    to_signed(17, 8),
    to_signed(-1, 8),
    to_signed(-25, 8),
    to_signed(-51, 8),
    to_signed(-73, 8),
    to_signed(-86, 8),
    to_signed(-86, 8),
    to_signed(-73, 8),
    to_signed(-50, 8),
    to_signed(-20, 8),
    to_signed(13, 8),
    to_signed(40, 8),
    to_signed(55, 8),
    to_signed(55, 8),
    to_signed(41, 8),
    to_signed(19, 8),
    to_signed(-2, 8),
    to_signed(-15, 8),
    to_signed(-17, 8),
    to_signed(-11, 8),
    to_signed(3, 8),
    to_signed(22, 8),
    to_signed(41, 8),
    to_signed(53, 8),
    to_signed(56, 8),
    to_signed(52, 8),
    to_signed(38, 8),
    to_signed(17, 8),
    to_signed(-4, 8),
    to_signed(-21, 8),
    to_signed(-35, 8),
    to_signed(-45, 8),
    to_signed(-51, 8),
    to_signed(-52, 8),
    to_signed(-50, 8),
    to_signed(-48, 8),
    to_signed(-45, 8),
    to_signed(-42, 8),
    to_signed(-39, 8),
    to_signed(-34, 8),
    to_signed(-26, 8),
    to_signed(-19, 8),
    to_signed(-17, 8),
    to_signed(-16, 8),
    to_signed(-13, 8),
    to_signed(-10, 8),
    to_signed(-7, 8),
    to_signed(-1, 8),
    to_signed(9, 8),
    to_signed(22, 8),
    to_signed(34, 8),
    to_signed(44, 8),
    to_signed(53, 8),
    to_signed(57, 8),
    to_signed(57, 8),
    to_signed(56, 8),
    to_signed(54, 8),
    to_signed(48, 8),
    to_signed(37, 8),
    to_signed(24, 8),
    to_signed(13, 8),
    to_signed(5, 8),
    to_signed(-1, 8),
    to_signed(-3, 8),
    to_signed(1, 8),
    to_signed(10, 8),
    to_signed(20, 8),
    to_signed(29, 8),
    to_signed(34, 8),
    to_signed(35, 8),
    to_signed(27, 8),
    to_signed(10, 8),
    to_signed(-16, 8),
    to_signed(-44, 8),
    to_signed(-69, 8),
    to_signed(-88, 8),
    to_signed(-95, 8),
    to_signed(-89, 8),
    to_signed(-70, 8),
    to_signed(-40, 8),
    to_signed(-7, 8),
    to_signed(24, 8),
    to_signed(45, 8),
    to_signed(50, 8),
    to_signed(40, 8),
    to_signed(22, 8),
    to_signed(2, 8),
    to_signed(-14, 8),
    to_signed(-22, 8),
    to_signed(-22, 8),
    to_signed(-13, 8),
    to_signed(3, 8),
    to_signed(21, 8),
    to_signed(35, 8),
    to_signed(43, 8),
    to_signed(44, 8),
    to_signed(37, 8),
    to_signed(24, 8),
    to_signed(6, 8),
    to_signed(-11, 8),
    to_signed(-24, 8),
    to_signed(-33, 8),
    to_signed(-41, 8),
    to_signed(-45, 8),
    to_signed(-47, 8),
    to_signed(-48, 8),
    to_signed(-48, 8),
    to_signed(-47, 8),
    to_signed(-46, 8),
    to_signed(-42, 8),
    to_signed(-35, 8),
    to_signed(-27, 8),
    to_signed(-20, 8),
    to_signed(-18, 8),
    to_signed(-17, 8),
    to_signed(-15, 8),
    to_signed(-14, 8),
    to_signed(-12, 8),
    to_signed(-5, 8),
    to_signed(8, 8),
    to_signed(21, 8),
    to_signed(32, 8),
    to_signed(41, 8),
    to_signed(49, 8),
    to_signed(54, 8),
    to_signed(58, 8),
    to_signed(60, 8),
    to_signed(56, 8),
    to_signed(46, 8),
    to_signed(33, 8),
    to_signed(23, 8),
    to_signed(16, 8),
    to_signed(10, 8),
    to_signed(4, 8),
    to_signed(5, 8),
    to_signed(12, 8),
    to_signed(22, 8),
    to_signed(32, 8),
    to_signed(39, 8),
    to_signed(41, 8),
    to_signed(36, 8),
    to_signed(24, 8),
    to_signed(4, 8),
    to_signed(-21, 8),
    to_signed(-47, 8),
    to_signed(-69, 8),
    to_signed(-84, 8),
    to_signed(-88, 8),
    to_signed(-77, 8),
    to_signed(-55, 8),
    to_signed(-26, 8),
    to_signed(4, 8),
    to_signed(29, 8),
    to_signed(42, 8),
    to_signed(42, 8),
    to_signed(31, 8),
    to_signed(17, 8),
    to_signed(2, 8),
    to_signed(-9, 8),
    to_signed(-12, 8),
    to_signed(-7, 8),
    to_signed(4, 8),
    to_signed(18, 8),
    to_signed(30, 8),
    to_signed(40, 8),
    to_signed(46, 8),
    to_signed(46, 8),
    to_signed(39, 8),
    to_signed(25, 8),
    to_signed(9, 8),
    to_signed(-4, 8),
    to_signed(-14, 8),
    to_signed(-23, 8),
    to_signed(-31, 8),
    to_signed(-37, 8),
    to_signed(-41, 8),
    to_signed(-46, 8),
    to_signed(-51, 8),
    to_signed(-52, 8),
    to_signed(-49, 8),
    to_signed(-42, 8),
    to_signed(-31, 8),
    to_signed(-20, 8),
    to_signed(-13, 8),
    to_signed(-13, 8),
    to_signed(-16, 8),
    to_signed(-17, 8),
    to_signed(-14, 8),
    to_signed(-7, 8),
    to_signed(5, 8),
    to_signed(21, 8),
    to_signed(37, 8),
    to_signed(49, 8),
    to_signed(56, 8),
    to_signed(60, 8),
    to_signed(60, 8),
    to_signed(57, 8),
    to_signed(51, 8),
    to_signed(41, 8),
    to_signed(29, 8),
    to_signed(18, 8),
    to_signed(11, 8),
    to_signed(4, 8),
    to_signed(0, 8),
    to_signed(0, 8),
    to_signed(5, 8),
    to_signed(12, 8),
    to_signed(18, 8),
    to_signed(23, 8),
    to_signed(26, 8),
    to_signed(26, 8),
    to_signed(21, 8),
    to_signed(11, 8),
    to_signed(-4, 8),
    to_signed(-25, 8),
    to_signed(-48, 8),
    to_signed(-68, 8),
    to_signed(-80, 8),
    to_signed(-81, 8),
    to_signed(-69, 8),
    to_signed(-48, 8),
    to_signed(-19, 8),
    to_signed(10, 8),
    to_signed(32, 8),
    to_signed(42, 8),
    to_signed(39, 8),
    to_signed(26, 8),
    to_signed(8, 8),
    to_signed(-9, 8),
    to_signed(-19, 8),
    to_signed(-19, 8),
    to_signed(-11, 8),
    to_signed(1, 8),
    to_signed(13, 8),
    to_signed(25, 8),
    to_signed(34, 8),
    to_signed(38, 8),
    to_signed(36, 8),
    to_signed(26, 8),
    to_signed(12, 8),
    to_signed(0, 8),
    to_signed(-10, 8),
    to_signed(-19, 8),
    to_signed(-28, 8),
    to_signed(-34, 8),
    to_signed(-37, 8),
    to_signed(-41, 8),
    to_signed(-47, 8),
    to_signed(-50, 8),
    to_signed(-48, 8),
    to_signed(-41, 8),
    to_signed(-32, 8),
    to_signed(-22, 8),
    to_signed(-13, 8),
    to_signed(-9, 8),
    to_signed(-12, 8),
    to_signed(-17, 8),
    to_signed(-18, 8),
    to_signed(-15, 8),
    to_signed(-8, 8),
    to_signed(6, 8),
    to_signed(24, 8),
    to_signed(40, 8),
    to_signed(50, 8),
    to_signed(54, 8),
    to_signed(54, 8),
    to_signed(51, 8),
    to_signed(46, 8),
    to_signed(39, 8),
    to_signed(30, 8),
    to_signed(22, 8),
    to_signed(16, 8),
    to_signed(14, 8),
    to_signed(14, 8),
    to_signed(15, 8),
    to_signed(18, 8),
    to_signed(22, 8),
    to_signed(26, 8),
    to_signed(29, 8),
    to_signed(34, 8),
    to_signed(38, 8),
    to_signed(39, 8),
    to_signed(35, 8),
    to_signed(25, 8),
    to_signed(7, 8),
    to_signed(-21, 8),
    to_signed(-51, 8),
    to_signed(-75, 8),
    to_signed(-86, 8),
    to_signed(-83, 8),
    to_signed(-68, 8),
    to_signed(-43, 8),
    to_signed(-11, 8),
    to_signed(18, 8),
    to_signed(37, 8),
    to_signed(42, 8),
    to_signed(34, 8),
    to_signed(19, 8),
    to_signed(3, 8),
    to_signed(-10, 8),
    to_signed(-14, 8),
    to_signed(-8, 8),
    to_signed(4, 8),
    to_signed(17, 8),
    to_signed(29, 8),
    to_signed(39, 8),
    to_signed(45, 8),
    to_signed(44, 8),
    to_signed(34, 8),
    to_signed(20, 8),
    to_signed(7, 8),
    to_signed(0, 8),
    to_signed(-6, 8),
    to_signed(-12, 8),
    to_signed(-19, 8),
    to_signed(-26, 8),
    to_signed(-33, 8),
    to_signed(-43, 8),
    to_signed(-53, 8),
    to_signed(-58, 8),
    to_signed(-56, 8),
    to_signed(-50, 8),
    to_signed(-42, 8),
    to_signed(-29, 8),
    to_signed(-17, 8),
    to_signed(-12, 8),
    to_signed(-15, 8),
    to_signed(-21, 8),
    to_signed(-23, 8),
    to_signed(-20, 8),
    to_signed(-10, 8),
    to_signed(7, 8),
    to_signed(26, 8),
    to_signed(40, 8),
    to_signed(49, 8),
    to_signed(56, 8),
    to_signed(59, 8),
    to_signed(57, 8),
    to_signed(51, 8),
    to_signed(42, 8),
    to_signed(34, 8),
    to_signed(28, 8),
    to_signed(23, 8),
    to_signed(18, 8),
    to_signed(14, 8),
    to_signed(13, 8),
    to_signed(16, 8),
    to_signed(23, 8),
    to_signed(28, 8),
    to_signed(31, 8),
    to_signed(32, 8),
    to_signed(29, 8),
    to_signed(20, 8),
    to_signed(7, 8),
    to_signed(-11, 8),
    to_signed(-37, 8),
    to_signed(-66, 8),
    to_signed(-89, 8),
    to_signed(-96, 8),
    to_signed(-91, 8),
    to_signed(-76, 8),
    to_signed(-53, 8),
    to_signed(-22, 8),
    to_signed(8, 8),
    to_signed(29, 8),
    to_signed(35, 8),
    to_signed(29, 8),
    to_signed(16, 8),
    to_signed(3, 8),
    to_signed(-7, 8),
    to_signed(-10, 8),
    to_signed(-6, 8),
    to_signed(5, 8),
    to_signed(18, 8),
    to_signed(30, 8),
    to_signed(39, 8),
    to_signed(42, 8),
    to_signed(37, 8),
    to_signed(25, 8),
    to_signed(9, 8),
    to_signed(-6, 8),
    to_signed(-16, 8),
    to_signed(-20, 8),
    to_signed(-24, 8),
    to_signed(-31, 8),
    to_signed(-39, 8),
    to_signed(-46, 8),
    to_signed(-51, 8),
    to_signed(-57, 8),
    to_signed(-61, 8),
    to_signed(-60, 8),
    to_signed(-54, 8),
    to_signed(-44, 8),
    to_signed(-33, 8),
    to_signed(-23, 8),
    to_signed(-18, 8),
    to_signed(-18, 8),
    to_signed(-20, 8),
    to_signed(-18, 8),
    to_signed(-12, 8),
    to_signed(-1, 8),
    to_signed(13, 8),
    to_signed(30, 8),
    to_signed(44, 8),
    to_signed(54, 8),
    to_signed(60, 8),
    to_signed(62, 8),
    to_signed(60, 8),
    to_signed(54, 8),
    to_signed(46, 8),
    to_signed(36, 8),
    to_signed(26, 8),
    to_signed(18, 8),
    to_signed(11, 8),
    to_signed(7, 8),
    to_signed(4, 8),
    to_signed(5, 8),
    to_signed(11, 8),
    to_signed(18, 8),
    to_signed(24, 8),
    to_signed(26, 8),
    to_signed(24, 8),
    to_signed(17, 8),
    to_signed(4, 8),
    to_signed(-13, 8),
    to_signed(-36, 8),
    to_signed(-61, 8),
    to_signed(-81, 8),
    to_signed(-89, 8),
    to_signed(-83, 8),
    to_signed(-68, 8),
    to_signed(-46, 8),
    to_signed(-17, 8),
    to_signed(13, 8),
    to_signed(34, 8),
    to_signed(39, 8),
    to_signed(31, 8),
    to_signed(17, 8),
    to_signed(1, 8),
    to_signed(-11, 8),
    to_signed(-16, 8),
    to_signed(-13, 8),
    to_signed(-5, 8),
    to_signed(6, 8),
    to_signed(18, 8),
    to_signed(29, 8),
    to_signed(35, 8),
    to_signed(33, 8),
    to_signed(28, 8),
    to_signed(19, 8),
    to_signed(10, 8),
    to_signed(-1, 8),
    to_signed(-9, 8),
    to_signed(-15, 8),
    to_signed(-21, 8),
    to_signed(-29, 8),
    to_signed(-37, 8),
    to_signed(-42, 8),
    to_signed(-46, 8),
    to_signed(-50, 8),
    to_signed(-52, 8),
    to_signed(-48, 8),
    to_signed(-39, 8),
    to_signed(-30, 8),
    to_signed(-23, 8),
    to_signed(-19, 8),
    to_signed(-17, 8),
    to_signed(-16, 8),
    to_signed(-15, 8),
    to_signed(-13, 8),
    to_signed(-8, 8),
    to_signed(1, 8),
    to_signed(15, 8),
    to_signed(31, 8),
    to_signed(44, 8),
    to_signed(50, 8),
    to_signed(53, 8),
    to_signed(51, 8),
    to_signed(48, 8),
    to_signed(43, 8),
    to_signed(38, 8),
    to_signed(33, 8),
    to_signed(29, 8),
    to_signed(27, 8),
    to_signed(26, 8),
    to_signed(22, 8),
    to_signed(17, 8),
    to_signed(16, 8),
    to_signed(21, 8),
    to_signed(29, 8),
    to_signed(35, 8),
    to_signed(38, 8),
    to_signed(37, 8),
    to_signed(30, 8),
    to_signed(17, 8),
    to_signed(-2, 8),
    to_signed(-27, 8),
    to_signed(-54, 8),
    to_signed(-75, 8),
    to_signed(-82, 8),
    to_signed(-76, 8),
    to_signed(-60, 8),
    to_signed(-38, 8),
    to_signed(-10, 8),
    to_signed(17, 8),
    to_signed(35, 8),
    to_signed(39, 8),
    to_signed(34, 8),
    to_signed(22, 8),
    to_signed(7, 8),
    to_signed(-8, 8),
    to_signed(-17, 8),
    to_signed(-17, 8),
    to_signed(-10, 8),
    to_signed(2, 8),
    to_signed(17, 8),
    to_signed(32, 8),
    to_signed(43, 8),
    to_signed(46, 8),
    to_signed(43, 8),
    to_signed(35, 8),
    to_signed(23, 8),
    to_signed(10, 8),
    to_signed(-2, 8),
    to_signed(-12, 8),
    to_signed(-22, 8),
    to_signed(-33, 8),
    to_signed(-43, 8),
    to_signed(-51, 8),
    to_signed(-57, 8),
    to_signed(-62, 8),
    to_signed(-64, 8),
    to_signed(-61, 8),
    to_signed(-52, 8),
    to_signed(-43, 8),
    to_signed(-37, 8),
    to_signed(-34, 8),
    to_signed(-33, 8),
    to_signed(-32, 8),
    to_signed(-29, 8),
    to_signed(-23, 8),
    to_signed(-14, 8),
    to_signed(-3, 8),
    to_signed(10, 8),
    to_signed(23, 8),
    to_signed(34, 8),
    to_signed(42, 8),
    to_signed(47, 8),
    to_signed(48, 8),
    to_signed(46, 8),
    to_signed(41, 8),
    to_signed(38, 8),
    to_signed(34, 8),
    to_signed(30, 8),
    to_signed(26, 8),
    to_signed(23, 8),
    to_signed(19, 8),
    to_signed(15, 8),
    to_signed(16, 8),
    to_signed(23, 8),
    to_signed(29, 8),
    to_signed(32, 8),
    to_signed(32, 8),
    to_signed(29, 8),
    to_signed(21, 8),
    to_signed(6, 8),
    to_signed(-17, 8),
    to_signed(-43, 8),
    to_signed(-68, 8),
    to_signed(-86, 8),
    to_signed(-91, 8),
    to_signed(-85, 8),
    to_signed(-71, 8),
    to_signed(-47, 8),
    to_signed(-17, 8),
    to_signed(13, 8),
    to_signed(32, 8),
    to_signed(37, 8),
    to_signed(33, 8),
    to_signed(21, 8),
    to_signed(7, 8),
    to_signed(-6, 8),
    to_signed(-16, 8),
    to_signed(-19, 8),
    to_signed(-14, 8),
    to_signed(-1, 8),
    to_signed(15, 8),
    to_signed(31, 8),
    to_signed(41, 8),
    to_signed(44, 8),
    to_signed(41, 8),
    to_signed(33, 8),
    to_signed(22, 8),
    to_signed(9, 8),
    to_signed(-6, 8),
    to_signed(-20, 8),
    to_signed(-32, 8),
    to_signed(-43, 8),
    to_signed(-51, 8),
    to_signed(-58, 8),
    to_signed(-62, 8),
    to_signed(-64, 8),
    to_signed(-62, 8),
    to_signed(-55, 8),
    to_signed(-45, 8),
    to_signed(-34, 8),
    to_signed(-25, 8),
    to_signed(-20, 8),
    to_signed(-16, 8),
    to_signed(-12, 8),
    to_signed(-7, 8),
    to_signed(-1, 8),
    to_signed(5, 8),
    to_signed(12, 8),
    to_signed(22, 8),
    to_signed(33, 8),
    to_signed(41, 8),
    to_signed(44, 8),
    to_signed(45, 8),
    to_signed(46, 8),
    to_signed(47, 8),
    to_signed(47, 8),
    to_signed(44, 8),
    to_signed(41, 8),
    to_signed(36, 8),
    to_signed(31, 8),
    to_signed(27, 8),
    to_signed(23, 8),
    to_signed(21, 8),
    to_signed(21, 8),
    to_signed(25, 8),
    to_signed(29, 8),
    to_signed(32, 8),
    to_signed(31, 8),
    to_signed(26, 8),
    to_signed(17, 8),
    to_signed(1, 8),
    to_signed(-20, 8),
    to_signed(-47, 8),
    to_signed(-73, 8),
    to_signed(-90, 8),
    to_signed(-93, 8),
    to_signed(-84, 8),
    to_signed(-68, 8),
    to_signed(-45, 8),
    to_signed(-17, 8),
    to_signed(10, 8),
    to_signed(26, 8),
    to_signed(29, 8),
    to_signed(24, 8),
    to_signed(13, 8),
    to_signed(1, 8),
    to_signed(-12, 8),
    to_signed(-19, 8),
    to_signed(-19, 8),
    to_signed(-11, 8),
    to_signed(2, 8),
    to_signed(16, 8),
    to_signed(29, 8),
    to_signed(40, 8),
    to_signed(45, 8),
    to_signed(44, 8),
    to_signed(39, 8),
    to_signed(31, 8),
    to_signed(20, 8),
    to_signed(6, 8),
    to_signed(-6, 8),
    to_signed(-16, 8),
    to_signed(-26, 8),
    to_signed(-38, 8),
    to_signed(-48, 8),
    to_signed(-53, 8),
    to_signed(-55, 8),
    to_signed(-54, 8),
    to_signed(-49, 8),
    to_signed(-40, 8),
    to_signed(-29, 8),
    to_signed(-21, 8),
    to_signed(-17, 8),
    to_signed(-15, 8),
    to_signed(-13, 8),
    to_signed(-10, 8),
    to_signed(-5, 8),
    to_signed(1, 8),
    to_signed(8, 8),
    to_signed(19, 8),
    to_signed(32, 8),
    to_signed(41, 8),
    to_signed(46, 8),
    to_signed(50, 8),
    to_signed(54, 8),
    to_signed(56, 8),
    to_signed(55, 8),
    to_signed(53, 8),
    to_signed(49, 8),
    to_signed(44, 8),
    to_signed(37, 8),
    to_signed(30, 8),
    to_signed(25, 8),
    to_signed(24, 8),
    to_signed(25, 8),
    to_signed(28, 8),
    to_signed(31, 8),
    to_signed(32, 8),
    to_signed(31, 8),
    to_signed(27, 8),
    to_signed(19, 8),
    to_signed(4, 8),
    to_signed(-18, 8),
    to_signed(-46, 8),
    to_signed(-72, 8),
    to_signed(-90, 8),
    to_signed(-96, 8),
    to_signed(-92, 8),
    to_signed(-80, 8),
    to_signed(-58, 8),
    to_signed(-27, 8),
    to_signed(5, 8),
    to_signed(26, 8),
    to_signed(33, 8),
    to_signed(29, 8),
    to_signed(20, 8),
    to_signed(8, 8),
    to_signed(-5, 8),
    to_signed(-14, 8),
    to_signed(-17, 8),
    to_signed(-14, 8),
    to_signed(-5, 8),
    to_signed(7, 8),
    to_signed(22, 8),
    to_signed(33, 8),
    to_signed(38, 8),
    to_signed(39, 8),
    to_signed(39, 8),
    to_signed(34, 8),
    to_signed(25, 8),
    to_signed(12, 8),
    to_signed(-1, 8),
    to_signed(-13, 8),
    to_signed(-26, 8),
    to_signed(-40, 8),
    to_signed(-51, 8),
    to_signed(-57, 8),
    to_signed(-58, 8),
    to_signed(-56, 8),
    to_signed(-49, 8),
    to_signed(-37, 8),
    to_signed(-25, 8),
    to_signed(-17, 8),
    to_signed(-13, 8),
    to_signed(-11, 8),
    to_signed(-10, 8),
    to_signed(-9, 8),
    to_signed(-7, 8),
    to_signed(-4, 8),
    to_signed(3, 8),
    to_signed(15, 8),
    to_signed(29, 8),
    to_signed(40, 8),
    to_signed(48, 8),
    to_signed(55, 8),
    to_signed(61, 8),
    to_signed(64, 8),
    to_signed(61, 8),
    to_signed(53, 8),
    to_signed(43, 8),
    to_signed(31, 8),
    to_signed(22, 8),
    to_signed(16, 8),
    to_signed(13, 8),
    to_signed(12, 8),
    to_signed(13, 8),
    to_signed(16, 8),
    to_signed(22, 8),
    to_signed(29, 8),
    to_signed(35, 8),
    to_signed(36, 8),
    to_signed(29, 8),
    to_signed(14, 8),
    to_signed(-7, 8),
    to_signed(-33, 8),
    to_signed(-59, 8),
    to_signed(-79, 8),
    to_signed(-87, 8),
    to_signed(-84, 8),
    to_signed(-71, 8),
    to_signed(-50, 8),
    to_signed(-20, 8),
    to_signed(11, 8),
    to_signed(32, 8),
    to_signed(40, 8),
    to_signed(38, 8),
    to_signed(30, 8),
    to_signed(17, 8),
    to_signed(1, 8),
    to_signed(-12, 8),
    to_signed(-21, 8),
    to_signed(-24, 8),
    to_signed(-18, 8),
    to_signed(-5, 8),
    to_signed(11, 8),
    to_signed(25, 8),
    to_signed(35, 8),
    to_signed(40, 8),
    to_signed(41, 8),
    to_signed(35, 8),
    to_signed(23, 8),
    to_signed(8, 8),
    to_signed(-5, 8),
    to_signed(-19, 8),
    to_signed(-35, 8),
    to_signed(-50, 8),
    to_signed(-59, 8),
    to_signed(-63, 8),
    to_signed(-63, 8),
    to_signed(-60, 8),
    to_signed(-53, 8),
    to_signed(-41, 8),
    to_signed(-30, 8),
    to_signed(-23, 8),
    to_signed(-19, 8),
    to_signed(-19, 8),
    to_signed(-20, 8),
    to_signed(-19, 8),
    to_signed(-15, 8),
    to_signed(-8, 8),
    to_signed(2, 8),
    to_signed(14, 8),
    to_signed(26, 8),
    to_signed(35, 8),
    to_signed(43, 8),
    to_signed(48, 8),
    to_signed(52, 8),
    to_signed(52, 8),
    to_signed(48, 8),
    to_signed(39, 8),
    to_signed(28, 8),
    to_signed(18, 8),
    to_signed(10, 8),
    to_signed(4, 8),
    to_signed(1, 8),
    to_signed(3, 8),
    to_signed(9, 8),
    to_signed(17, 8),
    to_signed(25, 8),
    to_signed(35, 8),
    to_signed(43, 8),
    to_signed(46, 8),
    to_signed(40, 8),
    to_signed(26, 8),
    to_signed(6, 8),
    to_signed(-20, 8),
    to_signed(-51, 8),
    to_signed(-78, 8),
    to_signed(-91, 8),
    to_signed(-87, 8),
    to_signed(-72, 8),
    to_signed(-51, 8),
    to_signed(-23, 8),
    to_signed(8, 8),
    to_signed(32, 8),
    to_signed(41, 8),
    to_signed(38, 8),
    to_signed(29, 8),
    to_signed(16, 8),
    to_signed(0, 8),
    to_signed(-14, 8),
    to_signed(-23, 8),
    to_signed(-24, 8),
    to_signed(-17, 8),
    to_signed(-3, 8),
    to_signed(14, 8),
    to_signed(30, 8),
    to_signed(43, 8),
    to_signed(49, 8),
    to_signed(47, 8),
    to_signed(39, 8),
    to_signed(24, 8),
    to_signed(8, 8),
    to_signed(-8, 8),
    to_signed(-23, 8),
    to_signed(-38, 8),
    to_signed(-50, 8),
    to_signed(-56, 8),
    to_signed(-57, 8),
    to_signed(-55, 8),
    to_signed(-52, 8),
    to_signed(-46, 8),
    to_signed(-38, 8),
    to_signed(-29, 8),
    to_signed(-24, 8),
    to_signed(-21, 8),
    to_signed(-20, 8),
    to_signed(-19, 8),
    to_signed(-18, 8),
    to_signed(-13, 8),
    to_signed(-4, 8),
    to_signed(6, 8),
    to_signed(18, 8),
    to_signed(28, 8),
    to_signed(35, 8),
    to_signed(39, 8),
    to_signed(41, 8),
    to_signed(43, 8),
    to_signed(42, 8),
    to_signed(37, 8),
    to_signed(27, 8),
    to_signed(17, 8),
    to_signed(8, 8),
    to_signed(0, 8),
    to_signed(-5, 8),
    to_signed(-5, 8),
    to_signed(-1, 8),
    to_signed(7, 8),
    to_signed(17, 8),
    to_signed(29, 8),
    to_signed(41, 8),
    to_signed(49, 8),
    to_signed(48, 8),
    to_signed(38, 8),
    to_signed(22, 8),
    to_signed(2, 8),
    to_signed(-24, 8),
    to_signed(-55, 8),
    to_signed(-83, 8),
    to_signed(-96, 8),
    to_signed(-92, 8),
    to_signed(-77, 8),
    to_signed(-54, 8),
    to_signed(-24, 8),
    to_signed(11, 8),
    to_signed(40, 8),
    to_signed(55, 8),
    to_signed(54, 8),
    to_signed(43, 8),
    to_signed(25, 8),
    to_signed(4, 8),
    to_signed(-14, 8),
    to_signed(-25, 8),
    to_signed(-28, 8),
    to_signed(-21, 8),
    to_signed(-6, 8),
    to_signed(13, 8),
    to_signed(33, 8),
    to_signed(49, 8),
    to_signed(57, 8),
    to_signed(55, 8),
    to_signed(44, 8),
    to_signed(29, 8),
    to_signed(13, 8),
    to_signed(-3, 8),
    to_signed(-19, 8),
    to_signed(-35, 8),
    to_signed(-47, 8),
    to_signed(-54, 8),
    to_signed(-53, 8),
    to_signed(-50, 8),
    to_signed(-45, 8),
    to_signed(-40, 8),
    to_signed(-32, 8),
    to_signed(-24, 8),
    to_signed(-18, 8),
    to_signed(-15, 8),
    to_signed(-13, 8),
    to_signed(-15, 8),
    to_signed(-19, 8),
    to_signed(-20, 8),
    to_signed(-14, 8),
    to_signed(-2, 8),
    to_signed(11, 8),
    to_signed(23, 8),
    to_signed(32, 8),
    to_signed(39, 8),
    to_signed(42, 8),
    to_signed(43, 8),
    to_signed(40, 8),
    to_signed(34, 8),
    to_signed(25, 8),
    to_signed(15, 8),
    to_signed(4, 8),
    to_signed(-2, 8),
    to_signed(-4, 8),
    to_signed(-2, 8),
    to_signed(4, 8),
    to_signed(14, 8),
    to_signed(25, 8),
    to_signed(37, 8),
    to_signed(47, 8),
    to_signed(55, 8),
    to_signed(54, 8),
    to_signed(45, 8),
    to_signed(28, 8),
    to_signed(4, 8),
    to_signed(-27, 8),
    to_signed(-61, 8),
    to_signed(-89, 8),
    to_signed(-101, 8),
    to_signed(-96, 8),
    to_signed(-81, 8),
    to_signed(-59, 8),
    to_signed(-28, 8),
    to_signed(9, 8),
    to_signed(43, 8),
    to_signed(64, 8),
    to_signed(68, 8),
    to_signed(57, 8),
    to_signed(35, 8),
    to_signed(10, 8),
    to_signed(-12, 8),
    to_signed(-27, 8),
    to_signed(-34, 8),
    to_signed(-30, 8),
    to_signed(-16, 8),
    to_signed(2, 8),
    to_signed(21, 8),
    to_signed(37, 8),
    to_signed(47, 8),
    to_signed(49, 8),
    to_signed(43, 8),
    to_signed(30, 8),
    to_signed(15, 8),
    to_signed(-1, 8),
    to_signed(-15, 8),
    to_signed(-27, 8),
    to_signed(-36, 8),
    to_signed(-41, 8),
    to_signed(-45, 8),
    to_signed(-47, 8),
    to_signed(-46, 8),
    to_signed(-41, 8),
    to_signed(-34, 8),
    to_signed(-29, 8),
    to_signed(-26, 8),
    to_signed(-26, 8),
    to_signed(-26, 8),
    to_signed(-25, 8),
    to_signed(-24, 8),
    to_signed(-21, 8),
    to_signed(-12, 8),
    to_signed(2, 8),
    to_signed(19, 8),
    to_signed(34, 8),
    to_signed(47, 8),
    to_signed(56, 8),
    to_signed(58, 8),
    to_signed(54, 8),
    to_signed(47, 8),
    to_signed(40, 8),
    to_signed(34, 8),
    to_signed(25, 8),
    to_signed(16, 8),
    to_signed(10, 8),
    to_signed(9, 8),
    to_signed(13, 8),
    to_signed(18, 8),
    to_signed(25, 8),
    to_signed(32, 8),
    to_signed(37, 8),
    to_signed(40, 8),
    to_signed(41, 8),
    to_signed(38, 8),
    to_signed(29, 8),
    to_signed(12, 8),
    to_signed(-11, 8),
    to_signed(-37, 8),
    to_signed(-65, 8),
    to_signed(-90, 8),
    to_signed(-102, 8),
    to_signed(-100, 8),
    to_signed(-87, 8),
    to_signed(-66, 8),
    to_signed(-36, 8),
    to_signed(0, 8),
    to_signed(32, 8),
    to_signed(51, 8),
    to_signed(53, 8),
    to_signed(41, 8),
    to_signed(19, 8),
    to_signed(-5, 8),
    to_signed(-24, 8),
    to_signed(-37, 8),
    to_signed(-40, 8),
    to_signed(-31, 8),
    to_signed(-12, 8),
    to_signed(10, 8),
    to_signed(31, 8),
    to_signed(46, 8),
    to_signed(53, 8),
    to_signed(50, 8),
    to_signed(37, 8),
    to_signed(20, 8),
    to_signed(4, 8),
    to_signed(-10, 8),
    to_signed(-23, 8),
    to_signed(-32, 8),
    to_signed(-37, 8),
    to_signed(-38, 8),
    to_signed(-40, 8),
    to_signed(-41, 8),
    to_signed(-39, 8),
    to_signed(-37, 8),
    to_signed(-37, 8),
    to_signed(-40, 8),
    to_signed(-41, 8),
    to_signed(-39, 8),
    to_signed(-36, 8),
    to_signed(-35, 8),
    to_signed(-33, 8),
    to_signed(-27, 8),
    to_signed(-14, 8),
    to_signed(3, 8),
    to_signed(22, 8),
    to_signed(40, 8),
    to_signed(53, 8),
    to_signed(60, 8),
    to_signed(60, 8),
    to_signed(57, 8),
    to_signed(50, 8),
    to_signed(42, 8),
    to_signed(32, 8),
    to_signed(22, 8),
    to_signed(12, 8),
    to_signed(6, 8),
    to_signed(6, 8),
    to_signed(10, 8),
    to_signed(15, 8),
    to_signed(21, 8),
    to_signed(27, 8),
    to_signed(32, 8),
    to_signed(35, 8),
    to_signed(37, 8),
    to_signed(37, 8),
    to_signed(31, 8),
    to_signed(17, 8),
    to_signed(-4, 8),
    to_signed(-30, 8),
    to_signed(-57, 8),
    to_signed(-83, 8),
    to_signed(-98, 8),
    to_signed(-100, 8),
    to_signed(-90, 8),
    to_signed(-70, 8),
    to_signed(-41, 8),
    to_signed(-4, 8),
    to_signed(30, 8),
    to_signed(49, 8),
    to_signed(51, 8),
    to_signed(42, 8),
    to_signed(23, 8),
    to_signed(-1, 8),
    to_signed(-21, 8),
    to_signed(-32, 8),
    to_signed(-35, 8),
    to_signed(-31, 8),
    to_signed(-17, 8),
    to_signed(5, 8),
    to_signed(29, 8),
    to_signed(46, 8),
    to_signed(53, 8),
    to_signed(51, 8),
    to_signed(42, 8),
    to_signed(25, 8),
    to_signed(7, 8),
    to_signed(-8, 8),
    to_signed(-21, 8),
    to_signed(-30, 8),
    to_signed(-34, 8),
    to_signed(-35, 8),
    to_signed(-36, 8),
    to_signed(-37, 8),
    to_signed(-36, 8),
    to_signed(-36, 8),
    to_signed(-36, 8),
    to_signed(-38, 8),
    to_signed(-38, 8),
    to_signed(-35, 8),
    to_signed(-32, 8),
    to_signed(-30, 8),
    to_signed(-26, 8),
    to_signed(-17, 8),
    to_signed(-4, 8),
    to_signed(10, 8),
    to_signed(24, 8),
    to_signed(37, 8),
    to_signed(49, 8),
    to_signed(57, 8),
    to_signed(60, 8),
    to_signed(59, 8),
    to_signed(52, 8),
    to_signed(41, 8),
    to_signed(30, 8),
    to_signed(20, 8),
    to_signed(10, 8),
    to_signed(2, 8),
    to_signed(0, 8),
    to_signed(6, 8),
    to_signed(13, 8),
    to_signed(19, 8),
    to_signed(27, 8),
    to_signed(37, 8),
    to_signed(43, 8),
    to_signed(45, 8),
    to_signed(45, 8),
    to_signed(43, 8),
    to_signed(36, 8),
    to_signed(21, 8),
    to_signed(0, 8),
    to_signed(-25, 8),
    to_signed(-52, 8),
    to_signed(-76, 8),
    to_signed(-90, 8),
    to_signed(-90, 8),
    to_signed(-76, 8),
    to_signed(-52, 8),
    to_signed(-21, 8),
    to_signed(10, 8),
    to_signed(34, 8),
    to_signed(49, 8),
    to_signed(52, 8),
    to_signed(42, 8),
    to_signed(21, 8),
    to_signed(-1, 8),
    to_signed(-16, 8),
    to_signed(-26, 8),
    to_signed(-29, 8),
    to_signed(-24, 8),
    to_signed(-9, 8),
    to_signed(11, 8),
    to_signed(27, 8),
    to_signed(37, 8),
    to_signed(42, 8),
    to_signed(41, 8),
    to_signed(31, 8),
    to_signed(18, 8),
    to_signed(5, 8),
    to_signed(-6, 8),
    to_signed(-15, 8),
    to_signed(-23, 8),
    to_signed(-27, 8),
    to_signed(-31, 8),
    to_signed(-34, 8),
    to_signed(-36, 8),
    to_signed(-35, 8),
    to_signed(-34, 8),
    to_signed(-35, 8),
    to_signed(-35, 8),
    to_signed(-33, 8),
    to_signed(-31, 8),
    to_signed(-31, 8),
    to_signed(-30, 8),
    to_signed(-25, 8),
    to_signed(-15, 8),
    to_signed(-2, 8),
    to_signed(8, 8),
    to_signed(19, 8),
    to_signed(32, 8),
    to_signed(41, 8),
    to_signed(46, 8),
    to_signed(47, 8),
    to_signed(45, 8),
    to_signed(39, 8),
    to_signed(33, 8),
    to_signed(26, 8),
    to_signed(19, 8),
    to_signed(11, 8),
    to_signed(7, 8),
    to_signed(8, 8),
    to_signed(11, 8),
    to_signed(13, 8),
    to_signed(16, 8),
    to_signed(21, 8),
    to_signed(25, 8),
    to_signed(26, 8),
    to_signed(27, 8),
    to_signed(28, 8),
    to_signed(27, 8),
    to_signed(20, 8),
    to_signed(6, 8),
    to_signed(-11, 8),
    to_signed(-33, 8),
    to_signed(-58, 8),
    to_signed(-80, 8),
    to_signed(-92, 8),
    to_signed(-90, 8),
    to_signed(-78, 8),
    to_signed(-58, 8),
    to_signed(-32, 8),
    to_signed(-4, 8),
    to_signed(23, 8),
    to_signed(42, 8),
    to_signed(46, 8),
    to_signed(36, 8),
    to_signed(19, 8),
    to_signed(1, 8),
    to_signed(-16, 8),
    to_signed(-30, 8),
    to_signed(-37, 8),
    to_signed(-33, 8),
    to_signed(-21, 8),
    to_signed(-8, 8),
    to_signed(4, 8),
    to_signed(15, 8),
    to_signed(23, 8),
    to_signed(26, 8),
    to_signed(21, 8),
    to_signed(14, 8),
    to_signed(6, 8),
    to_signed(-2, 8),
    to_signed(-9, 8),
    to_signed(-16, 8),
    to_signed(-22, 8),
    to_signed(-30, 8),
    to_signed(-37, 8),
    to_signed(-41, 8),
    to_signed(-42, 8),
    to_signed(-43, 8),
    to_signed(-43, 8),
    to_signed(-39, 8),
    to_signed(-33, 8),
    to_signed(-29, 8),
    to_signed(-27, 8),
    to_signed(-22, 8),
    to_signed(-14, 8),
    to_signed(-6, 8),
    to_signed(1, 8),
    to_signed(10, 8),
    to_signed(22, 8),
    to_signed(32, 8),
    to_signed(38, 8),
    to_signed(40, 8),
    to_signed(42, 8),
    to_signed(42, 8),
    to_signed(38, 8),
    to_signed(32, 8),
    to_signed(24, 8),
    to_signed(17, 8),
    to_signed(12, 8),
    to_signed(11, 8),
    to_signed(12, 8),
    to_signed(13, 8),
    to_signed(12, 8),
    to_signed(13, 8),
    to_signed(17, 8),
    to_signed(22, 8),
    to_signed(28, 8),
    to_signed(34, 8),
    to_signed(38, 8),
    to_signed(38, 8),
    to_signed(32, 8),
    to_signed(21, 8),
    to_signed(3, 8),
    to_signed(-22, 8),
    to_signed(-49, 8),
    to_signed(-70, 8),
    to_signed(-80, 8),
    to_signed(-78, 8),
    to_signed(-68, 8),
    to_signed(-50, 8),
    to_signed(-26, 8),
    to_signed(4, 8),
    to_signed(31, 8),
    to_signed(47, 8),
    to_signed(47, 8),
    to_signed(36, 8),
    to_signed(18, 8),
    to_signed(-4, 8),
    to_signed(-27, 8),
    to_signed(-46, 8),
    to_signed(-52, 8),
    to_signed(-46, 8),
    to_signed(-33, 8),
    to_signed(-17, 8),
    to_signed(0, 8),
    to_signed(18, 8),
    to_signed(32, 8),
    to_signed(38, 8),
    to_signed(38, 8),
    to_signed(35, 8),
    to_signed(31, 8),
    to_signed(23, 8),
    to_signed(10, 8),
    to_signed(-6, 8),
    to_signed(-21, 8),
    to_signed(-33, 8),
    to_signed(-42, 8),
    to_signed(-47, 8),
    to_signed(-46, 8),
    to_signed(-42, 8),
    to_signed(-36, 8),
    to_signed(-27, 8),
    to_signed(-19, 8),
    to_signed(-15, 8),
    to_signed(-13, 8),
    to_signed(-12, 8),
    to_signed(-11, 8),
    to_signed(-9, 8),
    to_signed(-3, 8),
    to_signed(8, 8),
    to_signed(20, 8),
    to_signed(31, 8),
    to_signed(42, 8),
    to_signed(50, 8),
    to_signed(51, 8),
    to_signed(47, 8),
    to_signed(41, 8),
    to_signed(33, 8),
    to_signed(24, 8),
    to_signed(15, 8),
    to_signed(8, 8),
    to_signed(5, 8),
    to_signed(3, 8),
    to_signed(3, 8),
    to_signed(7, 8),
    to_signed(16, 8),
    to_signed(25, 8),
    to_signed(34, 8),
    to_signed(42, 8),
    to_signed(51, 8),
    to_signed(57, 8),
    to_signed(54, 8),
    to_signed(44, 8),
    to_signed(26, 8),
    to_signed(1, 8),
    to_signed(-33, 8),
    to_signed(-65, 8),
    to_signed(-84, 8),
    to_signed(-91, 8),
    to_signed(-88, 8),
    to_signed(-75, 8),
    to_signed(-50, 8),
    to_signed(-16, 8),
    to_signed(18, 8),
    to_signed(42, 8),
    to_signed(51, 8),
    to_signed(47, 8),
    to_signed(34, 8),
    to_signed(13, 8),
    to_signed(-12, 8),
    to_signed(-33, 8),
    to_signed(-41, 8),
    to_signed(-36, 8),
    to_signed(-25, 8),
    to_signed(-12, 8),
    to_signed(2, 8),
    to_signed(18, 8),
    to_signed(33, 8),
    to_signed(41, 8),
    to_signed(43, 8),
    to_signed(38, 8),
    to_signed(30, 8),
    to_signed(19, 8),
    to_signed(6, 8),
    to_signed(-8, 8),
    to_signed(-22, 8),
    to_signed(-35, 8),
    to_signed(-47, 8),
    to_signed(-53, 8),
    to_signed(-52, 8),
    to_signed(-46, 8),
    to_signed(-39, 8),
    to_signed(-32, 8),
    to_signed(-24, 8),
    to_signed(-20, 8),
    to_signed(-20, 8),
    to_signed(-22, 8),
    to_signed(-23, 8),
    to_signed(-22, 8),
    to_signed(-18, 8),
    to_signed(-7, 8),
    to_signed(7, 8),
    to_signed(20, 8),
    to_signed(32, 8),
    to_signed(40, 8),
    to_signed(45, 8),
    to_signed(44, 8),
    to_signed(41, 8),
    to_signed(37, 8),
    to_signed(30, 8),
    to_signed(21, 8),
    to_signed(13, 8),
    to_signed(8, 8),
    to_signed(3, 8),
    to_signed(0, 8),
    to_signed(0, 8),
    to_signed(6, 8),
    to_signed(15, 8),
    to_signed(26, 8),
    to_signed(38, 8),
    to_signed(48, 8),
    to_signed(55, 8),
    to_signed(56, 8),
    to_signed(50, 8),
    to_signed(35, 8),
    to_signed(10, 8),
    to_signed(-25, 8),
    to_signed(-62, 8),
    to_signed(-88, 8),
    to_signed(-98, 8),
    to_signed(-95, 8),
    to_signed(-83, 8),
    to_signed(-59, 8),
    to_signed(-24, 8),
    to_signed(13, 8),
    to_signed(42, 8),
    to_signed(56, 8),
    to_signed(57, 8),
    to_signed(48, 8),
    to_signed(30, 8),
    to_signed(8, 8),
    to_signed(-12, 8),
    to_signed(-26, 8),
    to_signed(-30, 8),
    to_signed(-25, 8),
    to_signed(-15, 8),
    to_signed(-1, 8),
    to_signed(13, 8),
    to_signed(27, 8),
    to_signed(37, 8),
    to_signed(40, 8),
    to_signed(36, 8),
    to_signed(26, 8),
    to_signed(13, 8),
    to_signed(-1, 8),
    to_signed(-15, 8),
    to_signed(-26, 8),
    to_signed(-34, 8),
    to_signed(-39, 8),
    to_signed(-41, 8),
    to_signed(-41, 8),
    to_signed(-36, 8),
    to_signed(-29, 8),
    to_signed(-24, 8),
    to_signed(-20, 8),
    to_signed(-17, 8),
    to_signed(-16, 8),
    to_signed(-18, 8),
    to_signed(-19, 8),
    to_signed(-17, 8),
    to_signed(-12, 8),
    to_signed(-5, 8),
    to_signed(6, 8),
    to_signed(20, 8),
    to_signed(34, 8),
    to_signed(45, 8),
    to_signed(51, 8),
    to_signed(51, 8),
    to_signed(48, 8),
    to_signed(44, 8),
    to_signed(37, 8),
    to_signed(28, 8),
    to_signed(18, 8),
    to_signed(9, 8),
    to_signed(2, 8),
    to_signed(-2, 8),
    to_signed(-3, 8),
    to_signed(0, 8),
    to_signed(7, 8),
    to_signed(17, 8),
    to_signed(30, 8),
    to_signed(44, 8),
    to_signed(55, 8),
    to_signed(59, 8),
    to_signed(53, 8),
    to_signed(38, 8),
    to_signed(14, 8),
    to_signed(-19, 8),
    to_signed(-54, 8),
    to_signed(-81, 8),
    to_signed(-96, 8),
    to_signed(-97, 8),
    to_signed(-87, 8),
    to_signed(-67, 8),
    to_signed(-34, 8),
    to_signed(4, 8),
    to_signed(36, 8),
    to_signed(53, 8),
    to_signed(56, 8),
    to_signed(47, 8),
    to_signed(28, 8),
    to_signed(3, 8),
    to_signed(-20, 8),
    to_signed(-37, 8),
    to_signed(-45, 8),
    to_signed(-43, 8),
    to_signed(-32, 8),
    to_signed(-16, 8),
    to_signed(-1, 8),
    to_signed(14, 8),
    to_signed(26, 8),
    to_signed(32, 8),
    to_signed(28, 8),
    to_signed(18, 8),
    to_signed(5, 8),
    to_signed(-8, 8),
    to_signed(-18, 8),
    to_signed(-25, 8),
    to_signed(-31, 8),
    to_signed(-35, 8),
    to_signed(-37, 8),
    to_signed(-36, 8),
    to_signed(-32, 8),
    to_signed(-27, 8),
    to_signed(-24, 8),
    to_signed(-25, 8),
    to_signed(-26, 8),
    to_signed(-28, 8),
    to_signed(-30, 8),
    to_signed(-33, 8),
    to_signed(-31, 8),
    to_signed(-26, 8),
    to_signed(-17, 8),
    to_signed(-6, 8),
    to_signed(9, 8),
    to_signed(25, 8),
    to_signed(38, 8),
    to_signed(46, 8),
    to_signed(52, 8),
    to_signed(54, 8),
    to_signed(52, 8),
    to_signed(46, 8),
    to_signed(36, 8),
    to_signed(25, 8),
    to_signed(12, 8),
    to_signed(2, 8),
    to_signed(-4, 8),
    to_signed(-7, 8),
    to_signed(-5, 8),
    to_signed(2, 8),
    to_signed(13, 8),
    to_signed(26, 8),
    to_signed(38, 8),
    to_signed(49, 8),
    to_signed(54, 8),
    to_signed(50, 8),
    to_signed(36, 8),
    to_signed(12, 8),
    to_signed(-22, 8),
    to_signed(-60, 8),
    to_signed(-90, 8),
    to_signed(-104, 8),
    to_signed(-102, 8),
    to_signed(-91, 8),
    to_signed(-72, 8),
    to_signed(-43, 8),
    to_signed(-7, 8),
    to_signed(25, 8),
    to_signed(45, 8),
    to_signed(50, 8),
    to_signed(43, 8),
    to_signed(26, 8),
    to_signed(2, 8),
    to_signed(-20, 8),
    to_signed(-34, 8),
    to_signed(-38, 8),
    to_signed(-30, 8),
    to_signed(-11, 8),
    to_signed(14, 8),
    to_signed(34, 8),
    to_signed(45, 8),
    to_signed(49, 8),
    to_signed(48, 8),
    to_signed(38, 8),
    to_signed(22, 8),
    to_signed(5, 8),
    to_signed(-10, 8),
    to_signed(-20, 8),
    to_signed(-27, 8),
    to_signed(-29, 8),
    to_signed(-29, 8),
    to_signed(-27, 8),
    to_signed(-25, 8),
    to_signed(-21, 8),
    to_signed(-16, 8),
    to_signed(-15, 8),
    to_signed(-17, 8),
    to_signed(-22, 8),
    to_signed(-27, 8),
    to_signed(-30, 8),
    to_signed(-29, 8),
    to_signed(-21, 8),
    to_signed(-9, 8),
    to_signed(5, 8),
    to_signed(17, 8),
    to_signed(31, 8),
    to_signed(47, 8),
    to_signed(59, 8),
    to_signed(65, 8),
    to_signed(66, 8),
    to_signed(65, 8),
    to_signed(60, 8),
    to_signed(51, 8),
    to_signed(39, 8),
    to_signed(28, 8),
    to_signed(15, 8),
    to_signed(5, 8),
    to_signed(0, 8),
    to_signed(1, 8),
    to_signed(4, 8),
    to_signed(9, 8),
    to_signed(17, 8),
    to_signed(28, 8),
    to_signed(39, 8),
    to_signed(49, 8),
    to_signed(55, 8),
    to_signed(52, 8),
    to_signed(41, 8),
    to_signed(22, 8),
    to_signed(-5, 8),
    to_signed(-39, 8),
    to_signed(-71, 8),
    to_signed(-91, 8),
    to_signed(-94, 8),
    to_signed(-84, 8),
    to_signed(-67, 8),
    to_signed(-41, 8),
    to_signed(-8, 8),
    to_signed(23, 8),
    to_signed(43, 8),
    to_signed(49, 8),
    to_signed(43, 8),
    to_signed(27, 8),
    to_signed(5, 8),
    to_signed(-17, 8),
    to_signed(-33, 8),
    to_signed(-40, 8),
    to_signed(-38, 8),
    to_signed(-25, 8),
    to_signed(-4, 8),
    to_signed(19, 8),
    to_signed(33, 8),
    to_signed(39, 8),
    to_signed(39, 8),
    to_signed(32, 8),
    to_signed(18, 8),
    to_signed(2, 8),
    to_signed(-12, 8),
    to_signed(-20, 8),
    to_signed(-27, 8),
    to_signed(-32, 8),
    to_signed(-34, 8),
    to_signed(-34, 8),
    to_signed(-33, 8),
    to_signed(-31, 8),
    to_signed(-28, 8),
    to_signed(-27, 8),
    to_signed(-27, 8),
    to_signed(-28, 8),
    to_signed(-30, 8),
    to_signed(-33, 8),
    to_signed(-34, 8),
    to_signed(-30, 8),
    to_signed(-23, 8),
    to_signed(-13, 8),
    to_signed(-2, 8),
    to_signed(12, 8),
    to_signed(27, 8),
    to_signed(40, 8),
    to_signed(48, 8),
    to_signed(52, 8),
    to_signed(53, 8),
    to_signed(51, 8),
    to_signed(44, 8),
    to_signed(34, 8),
    to_signed(24, 8),
    to_signed(13, 8),
    to_signed(3, 8),
    to_signed(-4, 8),
    to_signed(-6, 8),
    to_signed(-3, 8),
    to_signed(2, 8),
    to_signed(10, 8),
    to_signed(20, 8),
    to_signed(31, 8),
    to_signed(41, 8),
    to_signed(49, 8),
    to_signed(51, 8),
    to_signed(44, 8),
    to_signed(27, 8),
    to_signed(1, 8),
    to_signed(-33, 8),
    to_signed(-70, 8),
    to_signed(-97, 8),
    to_signed(-105, 8),
    to_signed(-99, 8),
    to_signed(-85, 8),
    to_signed(-62, 8),
    to_signed(-29, 8),
    to_signed(6, 8),
    to_signed(33, 8),
    to_signed(46, 8),
    to_signed(45, 8),
    to_signed(32, 8),
    to_signed(12, 8),
    to_signed(-10, 8),
    to_signed(-27, 8),
    to_signed(-37, 8),
    to_signed(-38, 8),
    to_signed(-28, 8),
    to_signed(-7, 8),
    to_signed(18, 8),
    to_signed(37, 8),
    to_signed(46, 8),
    to_signed(46, 8),
    to_signed(42, 8),
    to_signed(31, 8),
    to_signed(16, 8),
    to_signed(0, 8),
    to_signed(-13, 8),
    to_signed(-21, 8),
    to_signed(-28, 8),
    to_signed(-31, 8),
    to_signed(-31, 8),
    to_signed(-29, 8),
    to_signed(-26, 8),
    to_signed(-22, 8),
    to_signed(-20, 8),
    to_signed(-19, 8),
    to_signed(-20, 8),
    to_signed(-24, 8),
    to_signed(-30, 8),
    to_signed(-33, 8),
    to_signed(-29, 8),
    to_signed(-21, 8),
    to_signed(-13, 8),
    to_signed(-4, 8),
    to_signed(10, 8),
    to_signed(26, 8),
    to_signed(41, 8),
    to_signed(51, 8),
    to_signed(56, 8),
    to_signed(56, 8),
    to_signed(50, 8),
    to_signed(42, 8),
    to_signed(34, 8),
    to_signed(24, 8),
    to_signed(14, 8),
    to_signed(5, 8),
    to_signed(-2, 8),
    to_signed(-5, 8),
    to_signed(-6, 8),
    to_signed(-3, 8),
    to_signed(3, 8),
    to_signed(13, 8),
    to_signed(26, 8),
    to_signed(37, 8),
    to_signed(46, 8),
    to_signed(48, 8),
    to_signed(43, 8),
    to_signed(31, 8),
    to_signed(14, 8),
    to_signed(-11, 8),
    to_signed(-43, 8),
    to_signed(-75, 8),
    to_signed(-95, 8),
    to_signed(-98, 8),
    to_signed(-91, 8),
    to_signed(-75, 8),
    to_signed(-50, 8),
    to_signed(-15, 8),
    to_signed(18, 8),
    to_signed(42, 8),
    to_signed(53, 8),
    to_signed(49, 8),
    to_signed(35, 8),
    to_signed(15, 8),
    to_signed(-5, 8),
    to_signed(-23, 8),
    to_signed(-35, 8),
    to_signed(-36, 8),
    to_signed(-25, 8),
    to_signed(-5, 8),
    to_signed(18, 8),
    to_signed(37, 8),
    to_signed(47, 8),
    to_signed(47, 8),
    to_signed(40, 8),
    to_signed(29, 8),
    to_signed(14, 8),
    to_signed(-1, 8),
    to_signed(-14, 8),
    to_signed(-24, 8),
    to_signed(-31, 8),
    to_signed(-33, 8),
    to_signed(-30, 8),
    to_signed(-25, 8),
    to_signed(-21, 8),
    to_signed(-18, 8),
    to_signed(-13, 8),
    to_signed(-9, 8),
    to_signed(-9, 8),
    to_signed(-13, 8),
    to_signed(-19, 8),
    to_signed(-22, 8),
    to_signed(-19, 8),
    to_signed(-13, 8),
    to_signed(-6, 8),
    to_signed(4, 8),
    to_signed(18, 8),
    to_signed(33, 8),
    to_signed(45, 8),
    to_signed(56, 8),
    to_signed(63, 8),
    to_signed(63, 8),
    to_signed(59, 8),
    to_signed(51, 8),
    to_signed(40, 8),
    to_signed(26, 8),
    to_signed(10, 8),
    to_signed(-1, 8),
    to_signed(-7, 8),
    to_signed(-7, 8),
    to_signed(-4, 8),
    to_signed(2, 8),
    to_signed(10, 8),
    to_signed(20, 8),
    to_signed(30, 8),
    to_signed(41, 8),
    to_signed(48, 8),
    to_signed(50, 8),
    to_signed(47, 8),
    to_signed(37, 8),
    to_signed(21, 8),
    to_signed(-4, 8),
    to_signed(-37, 8),
    to_signed(-68, 8),
    to_signed(-89, 8),
    to_signed(-95, 8),
    to_signed(-90, 8),
    to_signed(-73, 8),
    to_signed(-45, 8),
    to_signed(-9, 8),
    to_signed(23, 8),
    to_signed(44, 8),
    to_signed(50, 8),
    to_signed(44, 8),
    to_signed(29, 8),
    to_signed(8, 8),
    to_signed(-15, 8),
    to_signed(-34, 8),
    to_signed(-44, 8),
    to_signed(-43, 8),
    to_signed(-33, 8),
    to_signed(-16, 8),
    to_signed(3, 8),
    to_signed(18, 8),
    to_signed(24, 8),
    to_signed(22, 8),
    to_signed(17, 8),
    to_signed(10, 8),
    to_signed(1, 8),
    to_signed(-9, 8),
    to_signed(-19, 8),
    to_signed(-27, 8),
    to_signed(-32, 8),
    to_signed(-32, 8),
    to_signed(-28, 8),
    to_signed(-22, 8),
    to_signed(-18, 8),
    to_signed(-12, 8),
    to_signed(-5, 8),
    to_signed(0, 8),
    to_signed(-1, 8),
    to_signed(-7, 8),
    to_signed(-12, 8),
    to_signed(-17, 8),
    to_signed(-20, 8),
    to_signed(-21, 8),
    to_signed(-16, 8),
    to_signed(-5, 8),
    to_signed(9, 8),
    to_signed(26, 8),
    to_signed(42, 8),
    to_signed(56, 8),
    to_signed(61, 8),
    to_signed(58, 8),
    to_signed(51, 8),
    to_signed(43, 8),
    to_signed(33, 8),
    to_signed(19, 8),
    to_signed(4, 8),
    to_signed(-5, 8),
    to_signed(-9, 8),
    to_signed(-10, 8),
    to_signed(-8, 8),
    to_signed(-4, 8),
    to_signed(2, 8),
    to_signed(11, 8),
    to_signed(21, 8),
    to_signed(31, 8),
    to_signed(38, 8),
    to_signed(42, 8),
    to_signed(43, 8),
    to_signed(36, 8),
    to_signed(20, 8),
    to_signed(-5, 8),
    to_signed(-36, 8),
    to_signed(-66, 8),
    to_signed(-87, 8),
    to_signed(-95, 8),
    to_signed(-92, 8),
    to_signed(-78, 8),
    to_signed(-53, 8),
    to_signed(-19, 8),
    to_signed(13, 8),
    to_signed(35, 8),
    to_signed(43, 8),
    to_signed(42, 8),
    to_signed(30, 8),
    to_signed(8, 8),
    to_signed(-17, 8),
    to_signed(-35, 8),
    to_signed(-42, 8),
    to_signed(-40, 8),
    to_signed(-32, 8),
    to_signed(-19, 8),
    to_signed(-3, 8),
    to_signed(11, 8),
    to_signed(19, 8),
    to_signed(23, 8),
    to_signed(25, 8),
    to_signed(23, 8),
    to_signed(15, 8),
    to_signed(5, 8),
    to_signed(-3, 8),
    to_signed(-11, 8),
    to_signed(-18, 8),
    to_signed(-22, 8),
    to_signed(-22, 8),
    to_signed(-21, 8),
    to_signed(-21, 8),
    to_signed(-18, 8),
    to_signed(-13, 8),
    to_signed(-11, 8),
    to_signed(-13, 8),
    to_signed(-18, 8),
    to_signed(-23, 8),
    to_signed(-28, 8),
    to_signed(-30, 8),
    to_signed(-27, 8),
    to_signed(-17, 8),
    to_signed(-4, 8),
    to_signed(11, 8),
    to_signed(28, 8),
    to_signed(44, 8),
    to_signed(55, 8),
    to_signed(59, 8),
    to_signed(57, 8),
    to_signed(51, 8),
    to_signed(43, 8),
    to_signed(30, 8),
    to_signed(13, 8),
    to_signed(-3, 8),
    to_signed(-12, 8),
    to_signed(-16, 8),
    to_signed(-16, 8),
    to_signed(-15, 8),
    to_signed(-9, 8),
    to_signed(3, 8),
    to_signed(17, 8),
    to_signed(31, 8),
    to_signed(42, 8),
    to_signed(51, 8),
    to_signed(56, 8),
    to_signed(56, 8),
    to_signed(47, 8),
    to_signed(27, 8),
    to_signed(-2, 8),
    to_signed(-35, 8),
    to_signed(-68, 8),
    to_signed(-92, 8),
    to_signed(-102, 8),
    to_signed(-98, 8),
    to_signed(-81, 8),
    to_signed(-52, 8),
    to_signed(-14, 8),
    to_signed(20, 8),
    to_signed(43, 8),
    to_signed(55, 8),
    to_signed(53, 8),
    to_signed(35, 8),
    to_signed(5, 8),
    to_signed(-26, 8),
    to_signed(-47, 8),
    to_signed(-57, 8),
    to_signed(-57, 8),
    to_signed(-46, 8),
    to_signed(-24, 8),
    to_signed(1, 8),
    to_signed(21, 8),
    to_signed(34, 8),
    to_signed(39, 8),
    to_signed(38, 8),
    to_signed(30, 8),
    to_signed(18, 8),
    to_signed(6, 8),
    to_signed(-5, 8),
    to_signed(-15, 8),
    to_signed(-25, 8),
    to_signed(-30, 8),
    to_signed(-30, 8),
    to_signed(-29, 8),
    to_signed(-28, 8),
    to_signed(-22, 8),
    to_signed(-13, 8),
    to_signed(-8, 8),
    to_signed(-8, 8),
    to_signed(-12, 8),
    to_signed(-17, 8),
    to_signed(-23, 8),
    to_signed(-28, 8),
    to_signed(-26, 8),
    to_signed(-17, 8),
    to_signed(-3, 8),
    to_signed(15, 8),
    to_signed(36, 8),
    to_signed(54, 8),
    to_signed(65, 8),
    to_signed(70, 8),
    to_signed(70, 8),
    to_signed(64, 8),
    to_signed(51, 8),
    to_signed(31, 8),
    to_signed(10, 8),
    to_signed(-8, 8),
    to_signed(-17, 8),
    to_signed(-21, 8),
    to_signed(-20, 8),
    to_signed(-14, 8),
    to_signed(-3, 8),
    to_signed(10, 8),
    to_signed(24, 8),
    to_signed(36, 8),
    to_signed(45, 8),
    to_signed(52, 8),
    to_signed(56, 8),
    to_signed(55, 8),
    to_signed(44, 8),
    to_signed(23, 8),
    to_signed(-6, 8),
    to_signed(-39, 8),
    to_signed(-71, 8),
    to_signed(-94, 8),
    to_signed(-103, 8),
    to_signed(-96, 8),
    to_signed(-77, 8),
    to_signed(-48, 8),
    to_signed(-12, 8),
    to_signed(19, 8),
    to_signed(40, 8),
    to_signed(48, 8),
    to_signed(41, 8),
    to_signed(21, 8),
    to_signed(-6, 8),
    to_signed(-31, 8),
    to_signed(-50, 8),
    to_signed(-59, 8),
    to_signed(-58, 8),
    to_signed(-44, 8),
    to_signed(-24, 8),
    to_signed(-4, 8),
    to_signed(12, 8),
    to_signed(24, 8),
    to_signed(29, 8),
    to_signed(27, 8),
    to_signed(18, 8),
    to_signed(7, 8),
    to_signed(-3, 8),
    to_signed(-14, 8),
    to_signed(-24, 8),
    to_signed(-31, 8),
    to_signed(-33, 8),
    to_signed(-32, 8),
    to_signed(-31, 8),
    to_signed(-30, 8),
    to_signed(-24, 8),
    to_signed(-18, 8),
    to_signed(-15, 8),
    to_signed(-16, 8),
    to_signed(-18, 8),
    to_signed(-24, 8),
    to_signed(-32, 8),
    to_signed(-36, 8),
    to_signed(-33, 8),
    to_signed(-22, 8),
    to_signed(-6, 8),
    to_signed(14, 8),
    to_signed(36, 8),
    to_signed(54, 8),
    to_signed(64, 8),
    to_signed(69, 8),
    to_signed(68, 8),
    to_signed(60, 8),
    to_signed(45, 8),
    to_signed(27, 8),
    to_signed(10, 8),
    to_signed(-5, 8),
    to_signed(-14, 8),
    to_signed(-16, 8),
    to_signed(-12, 8),
    to_signed(-5, 8),
    to_signed(3, 8),
    to_signed(12, 8),
    to_signed(23, 8),
    to_signed(34, 8),
    to_signed(44, 8),
    to_signed(52, 8),
    to_signed(59, 8),
    to_signed(60, 8),
    to_signed(52, 8),
    to_signed(34, 8),
    to_signed(9, 8),
    to_signed(-21, 8),
    to_signed(-55, 8),
    to_signed(-82, 8),
    to_signed(-93, 8),
    to_signed(-89, 8),
    to_signed(-72, 8),
    to_signed(-44, 8),
    to_signed(-9, 8),
    to_signed(26, 8),
    to_signed(49, 8),
    to_signed(59, 8),
    to_signed(56, 8),
    to_signed(42, 8),
    to_signed(20, 8),
    to_signed(-4, 8),
    to_signed(-26, 8),
    to_signed(-41, 8),
    to_signed(-44, 8),
    to_signed(-36, 8),
    to_signed(-22, 8),
    to_signed(-6, 8),
    to_signed(10, 8),
    to_signed(22, 8),
    to_signed(27, 8),
    to_signed(24, 8),
    to_signed(18, 8),
    to_signed(12, 8),
    to_signed(6, 8),
    to_signed(-1, 8),
    to_signed(-9, 8),
    to_signed(-14, 8),
    to_signed(-17, 8),
    to_signed(-18, 8),
    to_signed(-19, 8),
    to_signed(-16, 8),
    to_signed(-11, 8),
    to_signed(-6, 8),
    to_signed(-5, 8),
    to_signed(-9, 8),
    to_signed(-15, 8),
    to_signed(-23, 8),
    to_signed(-28, 8),
    to_signed(-28, 8),
    to_signed(-23, 8),
    to_signed(-14, 8),
    to_signed(-1, 8),
    to_signed(18, 8),
    to_signed(36, 8),
    to_signed(48, 8),
    to_signed(55, 8),
    to_signed(60, 8),
    to_signed(60, 8),
    to_signed(52, 8),
    to_signed(38, 8),
    to_signed(23, 8),
    to_signed(9, 8),
    to_signed(-5, 8),
    to_signed(-13, 8),
    to_signed(-12, 8),
    to_signed(-7, 8),
    to_signed(-1, 8),
    to_signed(8, 8),
    to_signed(20, 8),
    to_signed(34, 8),
    to_signed(45, 8),
    to_signed(54, 8),
    to_signed(61, 8),
    to_signed(63, 8),
    to_signed(57, 8),
    to_signed(43, 8),
    to_signed(24, 8),
    to_signed(2, 8),
    to_signed(-26, 8),
    to_signed(-57, 8),
    to_signed(-80, 8),
    to_signed(-90, 8),
    to_signed(-88, 8),
    to_signed(-78, 8),
    to_signed(-58, 8),
    to_signed(-27, 8),
    to_signed(5, 8),
    to_signed(27, 8),
    to_signed(38, 8),
    to_signed(36, 8),
    to_signed(23, 8),
    to_signed(2, 8),
    to_signed(-22, 8),
    to_signed(-40, 8),
    to_signed(-50, 8),
    to_signed(-51, 8),
    to_signed(-43, 8),
    to_signed(-29, 8),
    to_signed(-11, 8),
    to_signed(7, 8),
    to_signed(19, 8),
    to_signed(24, 8),
    to_signed(23, 8),
    to_signed(21, 8),
    to_signed(17, 8),
    to_signed(9, 8),
    to_signed(-1, 8),
    to_signed(-9, 8),
    to_signed(-15, 8),
    to_signed(-18, 8),
    to_signed(-20, 8),
    to_signed(-20, 8),
    to_signed(-18, 8),
    to_signed(-15, 8),
    to_signed(-12, 8),
    to_signed(-11, 8),
    to_signed(-13, 8),
    to_signed(-18, 8),
    to_signed(-23, 8),
    to_signed(-26, 8),
    to_signed(-26, 8),
    to_signed(-24, 8),
    to_signed(-17, 8),
    to_signed(-4, 8),
    to_signed(12, 8),
    to_signed(27, 8),
    to_signed(39, 8),
    to_signed(50, 8),
    to_signed(59, 8),
    to_signed(59, 8),
    to_signed(52, 8),
    to_signed(43, 8),
    to_signed(33, 8),
    to_signed(20, 8),
    to_signed(5, 8),
    to_signed(-6, 8),
    to_signed(-9, 8),
    to_signed(-8, 8),
    to_signed(-4, 8),
    to_signed(5, 8),
    to_signed(17, 8),
    to_signed(29, 8),
    to_signed(39, 8),
    to_signed(46, 8),
    to_signed(50, 8),
    to_signed(48, 8),
    to_signed(39, 8),
    to_signed(28, 8),
    to_signed(13, 8),
    to_signed(-7, 8),
    to_signed(-35, 8),
    to_signed(-63, 8),
    to_signed(-82, 8),
    to_signed(-89, 8),
    to_signed(-86, 8),
    to_signed(-75, 8),
    to_signed(-51, 8),
    to_signed(-19, 8),
    to_signed(12, 8),
    to_signed(32, 8),
    to_signed(42, 8),
    to_signed(41, 8),
    to_signed(29, 8),
    to_signed(6, 8),
    to_signed(-19, 8),
    to_signed(-38, 8),
    to_signed(-48, 8),
    to_signed(-47, 8),
    to_signed(-36, 8),
    to_signed(-20, 8),
    to_signed(-1, 8),
    to_signed(16, 8),
    to_signed(28, 8),
    to_signed(33, 8),
    to_signed(32, 8),
    to_signed(27, 8),
    to_signed(19, 8),
    to_signed(8, 8),
    to_signed(-2, 8),
    to_signed(-13, 8),
    to_signed(-22, 8),
    to_signed(-26, 8),
    to_signed(-25, 8),
    to_signed(-20, 8),
    to_signed(-15, 8),
    to_signed(-7, 8),
    to_signed(0, 8),
    to_signed(2, 8),
    to_signed(-2, 8),
    to_signed(-11, 8),
    to_signed(-19, 8),
    to_signed(-25, 8),
    to_signed(-29, 8),
    to_signed(-27, 8),
    to_signed(-18, 8),
    to_signed(-4, 8),
    to_signed(11, 8),
    to_signed(26, 8),
    to_signed(41, 8),
    to_signed(52, 8),
    to_signed(59, 8),
    to_signed(59, 8),
    to_signed(53, 8),
    to_signed(45, 8),
    to_signed(32, 8),
    to_signed(16, 8),
    to_signed(0, 8),
    to_signed(-11, 8),
    to_signed(-17, 8),
    to_signed(-18, 8),
    to_signed(-15, 8),
    to_signed(-6, 8),
    to_signed(8, 8),
    to_signed(23, 8),
    to_signed(38, 8),
    to_signed(51, 8),
    to_signed(56, 8),
    to_signed(53, 8),
    to_signed(45, 8),
    to_signed(34, 8),
    to_signed(18, 8),
    to_signed(-2, 8),
    to_signed(-26, 8),
    to_signed(-47, 8),
    to_signed(-65, 8),
    to_signed(-77, 8),
    to_signed(-81, 8),
    to_signed(-73, 8),
    to_signed(-54, 8),
    to_signed(-28, 8),
    to_signed(-4, 8),
    to_signed(15, 8),
    to_signed(28, 8),
    to_signed(33, 8),
    to_signed(25, 8),
    to_signed(8, 8),
    to_signed(-10, 8),
    to_signed(-24, 8),
    to_signed(-35, 8),
    to_signed(-41, 8),
    to_signed(-39, 8),
    to_signed(-31, 8),
    to_signed(-17, 8),
    to_signed(0, 8),
    to_signed(16, 8),
    to_signed(28, 8),
    to_signed(32, 8),
    to_signed(32, 8),
    to_signed(28, 8),
    to_signed(22, 8),
    to_signed(14, 8),
    to_signed(7, 8),
    to_signed(1, 8),
    to_signed(-3, 8),
    to_signed(-7, 8),
    to_signed(-11, 8),
    to_signed(-12, 8),
    to_signed(-10, 8),
    to_signed(-6, 8),
    to_signed(-5, 8),
    to_signed(-6, 8),
    to_signed(-5, 8),
    to_signed(-7, 8),
    to_signed(-13, 8),
    to_signed(-19, 8),
    to_signed(-21, 8),
    to_signed(-16, 8),
    to_signed(-7, 8),
    to_signed(5, 8),
    to_signed(19, 8),
    to_signed(33, 8),
    to_signed(45, 8),
    to_signed(54, 8),
    to_signed(57, 8),
    to_signed(55, 8),
    to_signed(47, 8),
    to_signed(36, 8),
    to_signed(23, 8),
    to_signed(10, 8),
    to_signed(-2, 8),
    to_signed(-8, 8),
    to_signed(-10, 8),
    to_signed(-7, 8),
    to_signed(0, 8),
    to_signed(9, 8),
    to_signed(20, 8),
    to_signed(32, 8),
    to_signed(41, 8),
    to_signed(45, 8),
    to_signed(45, 8),
    to_signed(44, 8),
    to_signed(41, 8),
    to_signed(33, 8),
    to_signed(21, 8),
    to_signed(5, 8),
    to_signed(-15, 8),
    to_signed(-38, 8),
    to_signed(-62, 8),
    to_signed(-83, 8),
    to_signed(-94, 8),
    to_signed(-93, 8),
    to_signed(-79, 8),
    to_signed(-56, 8),
    to_signed(-29, 8),
    to_signed(-3, 8),
    to_signed(15, 8),
    to_signed(23, 8),
    to_signed(20, 8),
    to_signed(10, 8),
    to_signed(-9, 8),
    to_signed(-31, 8),
    to_signed(-50, 8),
    to_signed(-61, 8),
    to_signed(-63, 8),
    to_signed(-59, 8),
    to_signed(-46, 8),
    to_signed(-28, 8),
    to_signed(-9, 8),
    to_signed(6, 8),
    to_signed(17, 8),
    to_signed(24, 8),
    to_signed(24, 8),
    to_signed(19, 8),
    to_signed(10, 8),
    to_signed(-2, 8),
    to_signed(-14, 8),
    to_signed(-23, 8),
    to_signed(-27, 8),
    to_signed(-26, 8),
    to_signed(-23, 8),
    to_signed(-19, 8),
    to_signed(-16, 8),
    to_signed(-13, 8),
    to_signed(-13, 8),
    to_signed(-15, 8),
    to_signed(-20, 8),
    to_signed(-23, 8),
    to_signed(-24, 8),
    to_signed(-25, 8),
    to_signed(-22, 8),
    to_signed(-15, 8),
    to_signed(-3, 8),
    to_signed(10, 8),
    to_signed(22, 8),
    to_signed(31, 8),
    to_signed(36, 8),
    to_signed(36, 8),
    to_signed(32, 8),
    to_signed(26, 8),
    to_signed(19, 8),
    to_signed(9, 8),
    to_signed(-1, 8),
    to_signed(-8, 8),
    to_signed(-10, 8),
    to_signed(-6, 8),
    to_signed(1, 8),
    to_signed(10, 8),
    to_signed(19, 8),
    to_signed(27, 8),
    to_signed(32, 8),
    to_signed(37, 8),
    to_signed(42, 8),
    to_signed(47, 8),
    to_signed(49, 8),
    to_signed(46, 8),
    to_signed(39, 8),
    to_signed(28, 8),
    to_signed(13, 8),
    to_signed(-7, 8),
    to_signed(-29, 8),
    to_signed(-52, 8),
    to_signed(-72, 8),
    to_signed(-83, 8),
    to_signed(-84, 8),
    to_signed(-74, 8),
    to_signed(-56, 8),
    to_signed(-31, 8),
    to_signed(-3, 8),
    to_signed(20, 8),
    to_signed(32, 8),
    to_signed(32, 8),
    to_signed(22, 8),
    to_signed(5, 8),
    to_signed(-16, 8),
    to_signed(-37, 8),
    to_signed(-52, 8),
    to_signed(-59, 8),
    to_signed(-55, 8),
    to_signed(-44, 8),
    to_signed(-27, 8),
    to_signed(-8, 8),
    to_signed(11, 8),
    to_signed(25, 8),
    to_signed(33, 8),
    to_signed(36, 8),
    to_signed(34, 8),
    to_signed(30, 8),
    to_signed(21, 8),
    to_signed(10, 8),
    to_signed(0, 8),
    to_signed(-6, 8),
    to_signed(-9, 8),
    to_signed(-10, 8),
    to_signed(-11, 8),
    to_signed(-13, 8),
    to_signed(-15, 8),
    to_signed(-16, 8),
    to_signed(-17, 8),
    to_signed(-19, 8),
    to_signed(-23, 8),
    to_signed(-27, 8),
    to_signed(-26, 8),
    to_signed(-20, 8),
    to_signed(-9, 8),
    to_signed(3, 8),
    to_signed(16, 8),
    to_signed(27, 8),
    to_signed(37, 8),
    to_signed(42, 8),
    to_signed(45, 8),
    to_signed(44, 8),
    to_signed(40, 8),
    to_signed(32, 8),
    to_signed(25, 8),
    to_signed(20, 8),
    to_signed(17, 8),
    to_signed(17, 8),
    to_signed(20, 8),
    to_signed(25, 8),
    to_signed(30, 8),
    to_signed(32, 8),
    to_signed(32, 8),
    to_signed(32, 8),
    to_signed(35, 8),
    to_signed(41, 8),
    to_signed(47, 8),
    to_signed(51, 8),
    to_signed(51, 8),
    to_signed(45, 8),
    to_signed(30, 8),
    to_signed(8, 8),
    to_signed(-20, 8),
    to_signed(-50, 8),
    to_signed(-76, 8),
    to_signed(-92, 8),
    to_signed(-94, 8),
    to_signed(-86, 8),
    to_signed(-70, 8),
    to_signed(-44, 8),
    to_signed(-14, 8),
    to_signed(12, 8),
    to_signed(29, 8),
    to_signed(33, 8),
    to_signed(25, 8),
    to_signed(8, 8),
    to_signed(-13, 8),
    to_signed(-31, 8),
    to_signed(-42, 8),
    to_signed(-45, 8),
    to_signed(-41, 8),
    to_signed(-29, 8),
    to_signed(-11, 8),
    to_signed(7, 8),
    to_signed(21, 8),
    to_signed(28, 8),
    to_signed(31, 8),
    to_signed(30, 8),
    to_signed(27, 8),
    to_signed(20, 8),
    to_signed(14, 8),
    to_signed(10, 8),
    to_signed(6, 8),
    to_signed(2, 8),
    to_signed(-1, 8),
    to_signed(-5, 8),
    to_signed(-11, 8),
    to_signed(-17, 8),
    to_signed(-20, 8),
    to_signed(-21, 8),
    to_signed(-20, 8),
    to_signed(-18, 8),
    to_signed(-17, 8),
    to_signed(-16, 8),
    to_signed(-15, 8),
    to_signed(-10, 8),
    to_signed(0, 8),
    to_signed(11, 8),
    to_signed(22, 8),
    to_signed(32, 8),
    to_signed(41, 8),
    to_signed(48, 8),
    to_signed(52, 8),
    to_signed(52, 8),
    to_signed(47, 8),
    to_signed(39, 8),
    to_signed(31, 8),
    to_signed(24, 8),
    to_signed(17, 8),
    to_signed(12, 8),
    to_signed(9, 8),
    to_signed(8, 8),
    to_signed(11, 8),
    to_signed(15, 8),
    to_signed(18, 8),
    to_signed(22, 8),
    to_signed(27, 8),
    to_signed(35, 8),
    to_signed(44, 8),
    to_signed(51, 8),
    to_signed(53, 8),
    to_signed(49, 8),
    to_signed(36, 8),
    to_signed(17, 8),
    to_signed(-10, 8),
    to_signed(-43, 8),
    to_signed(-74, 8),
    to_signed(-92, 8),
    to_signed(-97, 8),
    to_signed(-90, 8),
    to_signed(-75, 8),
    to_signed(-49, 8),
    to_signed(-20, 8),
    to_signed(3, 8),
    to_signed(15, 8),
    to_signed(17, 8),
    to_signed(8, 8),
    to_signed(-9, 8),
    to_signed(-26, 8),
    to_signed(-39, 8),
    to_signed(-45, 8),
    to_signed(-45, 8),
    to_signed(-37, 8),
    to_signed(-23, 8),
    to_signed(-7, 8),
    to_signed(4, 8),
    to_signed(11, 8),
    to_signed(12, 8),
    to_signed(10, 8),
    to_signed(7, 8),
    to_signed(5, 8),
    to_signed(5, 8),
    to_signed(6, 8),
    to_signed(5, 8),
    to_signed(3, 8),
    to_signed(1, 8),
    to_signed(-1, 8),
    to_signed(-4, 8),
    to_signed(-9, 8),
    to_signed(-12, 8),
    to_signed(-12, 8),
    to_signed(-11, 8),
    to_signed(-11, 8),
    to_signed(-12, 8),
    to_signed(-13, 8),
    to_signed(-14, 8),
    to_signed(-15, 8),
    to_signed(-17, 8),
    to_signed(-16, 8),
    to_signed(-11, 8),
    to_signed(0, 8),
    to_signed(15, 8),
    to_signed(29, 8),
    to_signed(38, 8),
    to_signed(43, 8),
    to_signed(46, 8),
    to_signed(44, 8),
    to_signed(37, 8),
    to_signed(29, 8),
    to_signed(19, 8),
    to_signed(10, 8),
    to_signed(4, 8),
    to_signed(2, 8),
    to_signed(1, 8),
    to_signed(2, 8),
    to_signed(6, 8),
    to_signed(12, 8),
    to_signed(20, 8),
    to_signed(29, 8),
    to_signed(39, 8),
    to_signed(49, 8),
    to_signed(56, 8),
    to_signed(57, 8),
    to_signed(51, 8),
    to_signed(36, 8),
    to_signed(12, 8),
    to_signed(-19, 8),
    to_signed(-52, 8),
    to_signed(-80, 8),
    to_signed(-96, 8),
    to_signed(-98, 8),
    to_signed(-87, 8),
    to_signed(-63, 8),
    to_signed(-32, 8),
    to_signed(-2, 8),
    to_signed(20, 8),
    to_signed(28, 8),
    to_signed(24, 8),
    to_signed(9, 8),
    to_signed(-15, 8),
    to_signed(-38, 8),
    to_signed(-55, 8),
    to_signed(-64, 8),
    to_signed(-63, 8),
    to_signed(-50, 8),
    to_signed(-29, 8),
    to_signed(-5, 8),
    to_signed(15, 8),
    to_signed(27, 8),
    to_signed(29, 8),
    to_signed(23, 8),
    to_signed(15, 8),
    to_signed(7, 8),
    to_signed(1, 8),
    to_signed(-4, 8),
    to_signed(-8, 8),
    to_signed(-12, 8),
    to_signed(-13, 8),
    to_signed(-11, 8),
    to_signed(-8, 8),
    to_signed(-5, 8),
    to_signed(-3, 8),
    to_signed(-1, 8),
    to_signed(1, 8),
    to_signed(-1, 8),
    to_signed(-3, 8),
    to_signed(-4, 8),
    to_signed(-6, 8),
    to_signed(-11, 8),
    to_signed(-13, 8),
    to_signed(-12, 8),
    to_signed(-7, 8),
    to_signed(-1, 8),
    to_signed(9, 8),
    to_signed(22, 8),
    to_signed(36, 8),
    to_signed(47, 8),
    to_signed(52, 8),
    to_signed(51, 8),
    to_signed(45, 8),
    to_signed(37, 8),
    to_signed(30, 8),
    to_signed(21, 8),
    to_signed(12, 8),
    to_signed(4, 8),
    to_signed(0, 8),
    to_signed(0, 8),
    to_signed(3, 8),
    to_signed(9, 8),
    to_signed(18, 8),
    to_signed(31, 8),
    to_signed(43, 8),
    to_signed(49, 8),
    to_signed(48, 8),
    to_signed(43, 8),
    to_signed(35, 8),
    to_signed(23, 8),
    to_signed(3, 8),
    to_signed(-22, 8),
    to_signed(-50, 8),
    to_signed(-74, 8),
    to_signed(-87, 8),
    to_signed(-87, 8),
    to_signed(-76, 8),
    to_signed(-55, 8),
    to_signed(-27, 8),
    to_signed(1, 8),
    to_signed(22, 8),
    to_signed(30, 8),
    to_signed(26, 8),
    to_signed(10, 8),
    to_signed(-13, 8),
    to_signed(-38, 8),
    to_signed(-59, 8),
    to_signed(-70, 8),
    to_signed(-70, 8),
    to_signed(-57, 8),
    to_signed(-36, 8),
    to_signed(-13, 8),
    to_signed(7, 8),
    to_signed(20, 8),
    to_signed(25, 8),
    to_signed(22, 8),
    to_signed(16, 8),
    to_signed(9, 8),
    to_signed(4, 8),
    to_signed(0, 8),
    to_signed(-3, 8),
    to_signed(-5, 8),
    to_signed(-7, 8),
    to_signed(-9, 8),
    to_signed(-10, 8),
    to_signed(-10, 8),
    to_signed(-7, 8),
    to_signed(-2, 8),
    to_signed(2, 8),
    to_signed(3, 8),
    to_signed(1, 8),
    to_signed(0, 8),
    to_signed(-4, 8),
    to_signed(-8, 8),
    to_signed(-11, 8),
    to_signed(-11, 8),
    to_signed(-7, 8),
    to_signed(0, 8),
    to_signed(9, 8),
    to_signed(21, 8),
    to_signed(34, 8),
    to_signed(45, 8),
    to_signed(53, 8),
    to_signed(53, 8),
    to_signed(49, 8),
    to_signed(42, 8),
    to_signed(35, 8),
    to_signed(28, 8),
    to_signed(20, 8),
    to_signed(12, 8),
    to_signed(4, 8),
    to_signed(-2, 8),
    to_signed(-5, 8),
    to_signed(-3, 8),
    to_signed(6, 8),
    to_signed(21, 8),
    to_signed(38, 8),
    to_signed(51, 8),
    to_signed(60, 8),
    to_signed(63, 8),
    to_signed(60, 8),
    to_signed(47, 8),
    to_signed(26, 8),
    to_signed(-2, 8),
    to_signed(-33, 8),
    to_signed(-62, 8),
    to_signed(-83, 8),
    to_signed(-89, 8),
    to_signed(-83, 8),
    to_signed(-66, 8),
    to_signed(-41, 8),
    to_signed(-13, 8),
    to_signed(11, 8),
    to_signed(24, 8),
    to_signed(26, 8),
    to_signed(16, 8),
    to_signed(0, 8),
    to_signed(-18, 8),
    to_signed(-34, 8),
    to_signed(-48, 8),
    to_signed(-57, 8),
    to_signed(-57, 8),
    to_signed(-47, 8),
    to_signed(-31, 8),
    to_signed(-14, 8),
    to_signed(1, 8),
    to_signed(13, 8),
    to_signed(22, 8),
    to_signed(26, 8),
    to_signed(24, 8),
    to_signed(19, 8),
    to_signed(13, 8),
    to_signed(8, 8),
    to_signed(2, 8),
    to_signed(-4, 8),
    to_signed(-10, 8),
    to_signed(-14, 8),
    to_signed(-15, 8),
    to_signed(-12, 8),
    to_signed(-5, 8),
    to_signed(1, 8),
    to_signed(4, 8),
    to_signed(4, 8),
    to_signed(3, 8),
    to_signed(-1, 8),
    to_signed(-8, 8),
    to_signed(-13, 8),
    to_signed(-15, 8),
    to_signed(-12, 8),
    to_signed(-5, 8),
    to_signed(6, 8),
    to_signed(17, 8),
    to_signed(27, 8),
    to_signed(36, 8),
    to_signed(44, 8),
    to_signed(47, 8),
    to_signed(46, 8),
    to_signed(41, 8),
    to_signed(33, 8),
    to_signed(21, 8),
    to_signed(10, 8),
    to_signed(1, 8),
    to_signed(-6, 8),
    to_signed(-12, 8),
    to_signed(-13, 8),
    to_signed(-9, 8),
    to_signed(1, 8),
    to_signed(15, 8),
    to_signed(28, 8),
    to_signed(39, 8),
    to_signed(46, 8),
    to_signed(49, 8),
    to_signed(48, 8),
    to_signed(41, 8),
    to_signed(28, 8),
    to_signed(10, 8),
    to_signed(-8, 8),
    to_signed(-26, 8),
    to_signed(-42, 8),
    to_signed(-58, 8),
    to_signed(-73, 8),
    to_signed(-82, 8),
    to_signed(-83, 8),
    to_signed(-77, 8),
    to_signed(-64, 8),
    to_signed(-45, 8),
    to_signed(-22, 8),
    to_signed(-3, 8),
    to_signed(9, 8),
    to_signed(15, 8),
    to_signed(12, 8),
    to_signed(0, 8),
    to_signed(-16, 8),
    to_signed(-32, 8),
    to_signed(-47, 8),
    to_signed(-58, 8),
    to_signed(-62, 8),
    to_signed(-56, 8),
    to_signed(-42, 8),
    to_signed(-21, 8),
    to_signed(1, 8),
    to_signed(19, 8),
    to_signed(29, 8),
    to_signed(31, 8),
    to_signed(24, 8),
    to_signed(12, 8),
    to_signed(-1, 8),
    to_signed(-10, 8),
    to_signed(-16, 8),
    to_signed(-18, 8),
    to_signed(-17, 8),
    to_signed(-12, 8),
    to_signed(-6, 8),
    to_signed(0, 8),
    to_signed(4, 8),
    to_signed(7, 8),
    to_signed(6, 8),
    to_signed(1, 8),
    to_signed(-4, 8),
    to_signed(-8, 8),
    to_signed(-10, 8),
    to_signed(-11, 8),
    to_signed(-9, 8),
    to_signed(-4, 8),
    to_signed(5, 8),
    to_signed(14, 8),
    to_signed(22, 8),
    to_signed(28, 8),
    to_signed(33, 8),
    to_signed(37, 8),
    to_signed(36, 8),
    to_signed(33, 8),
    to_signed(29, 8),
    to_signed(23, 8),
    to_signed(16, 8),
    to_signed(10, 8),
    to_signed(7, 8),
    to_signed(7, 8),
    to_signed(7, 8),
    to_signed(11, 8),
    to_signed(17, 8),
    to_signed(23, 8),
    to_signed(28, 8),
    to_signed(34, 8),
    to_signed(40, 8),
    to_signed(42, 8),
    to_signed(41, 8),
    to_signed(37, 8),
    to_signed(29, 8),
    to_signed(18, 8),
    to_signed(5, 8),
    to_signed(-10, 8),
    to_signed(-27, 8),
    to_signed(-46, 8),
    to_signed(-64, 8),
    to_signed(-75, 8),
    to_signed(-77, 8),
    to_signed(-68, 8),
    to_signed(-51, 8),
    to_signed(-30, 8),
    to_signed(-8, 8),
    to_signed(11, 8),
    to_signed(23, 8),
    to_signed(23, 8),
    to_signed(14, 8),
    to_signed(-1, 8),
    to_signed(-19, 8),
    to_signed(-38, 8),
    to_signed(-55, 8),
    to_signed(-62, 8),
    to_signed(-58, 8),
    to_signed(-45, 8),
    to_signed(-28, 8),
    to_signed(-11, 8),
    to_signed(4, 8),
    to_signed(17, 8),
    to_signed(24, 8),
    to_signed(24, 8),
    to_signed(20, 8),
    to_signed(15, 8),
    to_signed(8, 8),
    to_signed(2, 8),
    to_signed(-1, 8),
    to_signed(-2, 8),
    to_signed(-3, 8),
    to_signed(-5, 8),
    to_signed(-7, 8),
    to_signed(-9, 8),
    to_signed(-13, 8),
    to_signed(-15, 8),
    to_signed(-15, 8),
    to_signed(-15, 8),
    to_signed(-15, 8),
    to_signed(-15, 8),
    to_signed(-15, 8),
    to_signed(-12, 8),
    to_signed(-7, 8),
    to_signed(1, 8),
    to_signed(12, 8),
    to_signed(23, 8),
    to_signed(33, 8),
    to_signed(38, 8),
    to_signed(40, 8),
    to_signed(40, 8),
    to_signed(37, 8),
    to_signed(29, 8),
    to_signed(20, 8),
    to_signed(11, 8),
    to_signed(6, 8),
    to_signed(2, 8),
    to_signed(0, 8),
    to_signed(3, 8),
    to_signed(10, 8),
    to_signed(18, 8),
    to_signed(25, 8),
    to_signed(30, 8),
    to_signed(34, 8),
    to_signed(36, 8),
    to_signed(37, 8),
    to_signed(37, 8),
    to_signed(36, 8),
    to_signed(33, 8),
    to_signed(27, 8),
    to_signed(15, 8),
    to_signed(-2, 8),
    to_signed(-23, 8),
    to_signed(-44, 8),
    to_signed(-63, 8),
    to_signed(-75, 8),
    to_signed(-77, 8),
    to_signed(-70, 8),
    to_signed(-53, 8),
    to_signed(-30, 8),
    to_signed(-5, 8),
    to_signed(15, 8),
    to_signed(27, 8),
    to_signed(28, 8),
    to_signed(18, 8),
    to_signed(-3, 8),
    to_signed(-27, 8),
    to_signed(-47, 8),
    to_signed(-57, 8),
    to_signed(-57, 8),
    to_signed(-48, 8),
    to_signed(-31, 8),
    to_signed(-12, 8),
    to_signed(7, 8),
    to_signed(20, 8),
    to_signed(27, 8),
    to_signed(28, 8),
    to_signed(26, 8),
    to_signed(20, 8),
    to_signed(11, 8),
    to_signed(4, 8),
    to_signed(1, 8),
    to_signed(2, 8),
    to_signed(2, 8),
    to_signed(2, 8),
    to_signed(1, 8),
    to_signed(0, 8),
    to_signed(0, 8),
    to_signed(0, 8),
    to_signed(2, 8),
    to_signed(3, 8),
    to_signed(4, 8),
    to_signed(2, 8),
    to_signed(-1, 8),
    to_signed(-3, 8),
    to_signed(-2, 8),
    to_signed(2, 8),
    to_signed(9, 8),
    to_signed(19, 8),
    to_signed(31, 8),
    to_signed(42, 8),
    to_signed(49, 8),
    to_signed(52, 8),
    to_signed(51, 8),
    to_signed(47, 8),
    to_signed(38, 8),
    to_signed(27, 8),
    to_signed(14, 8),
    to_signed(3, 8),
    to_signed(-5, 8),
    to_signed(-7, 8),
    to_signed(-5, 8),
    to_signed(1, 8),
    to_signed(11, 8),
    to_signed(25, 8),
    to_signed(37, 8),
    to_signed(45, 8),
    to_signed(51, 8),
    to_signed(55, 8),
    to_signed(54, 8),
    to_signed(49, 8),
    to_signed(39, 8),
    to_signed(23, 8),
    to_signed(2, 8),
    to_signed(-25, 8),
    to_signed(-53, 8),
    to_signed(-77, 8),
    to_signed(-92, 8),
    to_signed(-93, 8),
    to_signed(-81, 8),
    to_signed(-57, 8),
    to_signed(-26, 8),
    to_signed(5, 8),
    to_signed(27, 8),
    to_signed(37, 8),
    to_signed(32, 8),
    to_signed(16, 8),
    to_signed(-6, 8),
    to_signed(-30, 8),
    to_signed(-50, 8),
    to_signed(-62, 8),
    to_signed(-61, 8),
    to_signed(-47, 8),
    to_signed(-25, 8),
    to_signed(-1, 8),
    to_signed(21, 8),
    to_signed(36, 8),
    to_signed(40, 8),
    to_signed(34, 8),
    to_signed(21, 8),
    to_signed(7, 8),
    to_signed(-7, 8),
    to_signed(-16, 8),
    to_signed(-20, 8),
    to_signed(-20, 8),
    to_signed(-18, 8),
    to_signed(-15, 8),
    to_signed(-10, 8),
    to_signed(-5, 8),
    to_signed(-1, 8),
    to_signed(1, 8),
    to_signed(1, 8),
    to_signed(-1, 8),
    to_signed(-5, 8),
    to_signed(-10, 8),
    to_signed(-15, 8),
    to_signed(-20, 8),
    to_signed(-21, 8),
    to_signed(-18, 8),
    to_signed(-10, 8),
    to_signed(2, 8),
    to_signed(17, 8),
    to_signed(32, 8),
    to_signed(47, 8),
    to_signed(56, 8),
    to_signed(58, 8),
    to_signed(51, 8),
    to_signed(40, 8),
    to_signed(28, 8),
    to_signed(16, 8),
    to_signed(5, 8),
    to_signed(-5, 8),
    to_signed(-11, 8),
    to_signed(-10, 8),
    to_signed(-2, 8),
    to_signed(11, 8),
    to_signed(24, 8),
    to_signed(34, 8),
    to_signed(42, 8),
    to_signed(47, 8),
    to_signed(47, 8),
    to_signed(41, 8),
    to_signed(30, 8),
    to_signed(17, 8),
    to_signed(2, 8),
    to_signed(-16, 8),
    to_signed(-35, 8),
    to_signed(-55, 8),
    to_signed(-73, 8),
    to_signed(-84, 8),
    to_signed(-88, 8),
    to_signed(-81, 8),
    to_signed(-61, 8),
    to_signed(-33, 8),
    to_signed(-4, 8),
    to_signed(17, 8),
    to_signed(27, 8),
    to_signed(25, 8),
    to_signed(14, 8),
    to_signed(-5, 8),
    to_signed(-26, 8),
    to_signed(-44, 8),
    to_signed(-54, 8),
    to_signed(-53, 8),
    to_signed(-44, 8),
    to_signed(-29, 8),
    to_signed(-12, 8),
    to_signed(6, 8),
    to_signed(20, 8),
    to_signed(24, 8),
    to_signed(20, 8),
    to_signed(12, 8),
    to_signed(4, 8),
    to_signed(-5, 8),
    to_signed(-12, 8),
    to_signed(-15, 8),
    to_signed(-16, 8),
    to_signed(-14, 8),
    to_signed(-13, 8),
    to_signed(-10, 8),
    to_signed(-6, 8),
    to_signed(0, 8),
    to_signed(4, 8),
    to_signed(4, 8),
    to_signed(3, 8),
    to_signed(2, 8),
    to_signed(-1, 8),
    to_signed(-7, 8),
    to_signed(-14, 8),
    to_signed(-19, 8),
    to_signed(-21, 8),
    to_signed(-15, 8),
    to_signed(-4, 8),
    to_signed(13, 8),
    to_signed(31, 8),
    to_signed(48, 8),
    to_signed(59, 8),
    to_signed(63, 8),
    to_signed(59, 8),
    to_signed(50, 8),
    to_signed(40, 8),
    to_signed(30, 8),
    to_signed(19, 8),
    to_signed(9, 8),
    to_signed(2, 8),
    to_signed(0, 8),
    to_signed(3, 8),
    to_signed(12, 8),
    to_signed(23, 8),
    to_signed(32, 8),
    to_signed(37, 8),
    to_signed(39, 8),
    to_signed(40, 8),
    to_signed(39, 8),
    to_signed(34, 8),
    to_signed(24, 8),
    to_signed(10, 8),
    to_signed(-7, 8),
    to_signed(-26, 8),
    to_signed(-46, 8),
    to_signed(-66, 8),
    to_signed(-82, 8),
    to_signed(-89, 8),
    to_signed(-83, 8),
    to_signed(-65, 8),
    to_signed(-41, 8),
    to_signed(-15, 8),
    to_signed(7, 8),
    to_signed(20, 8),
    to_signed(19, 8),
    to_signed(7, 8),
    to_signed(-13, 8),
    to_signed(-35, 8),
    to_signed(-54, 8),
    to_signed(-66, 8),
    to_signed(-66, 8),
    to_signed(-55, 8),
    to_signed(-37, 8),
    to_signed(-14, 8),
    to_signed(9, 8),
    to_signed(23, 8),
    to_signed(28, 8),
    to_signed(26, 8),
    to_signed(19, 8),
    to_signed(9, 8),
    to_signed(-1, 8),
    to_signed(-8, 8),
    to_signed(-13, 8),
    to_signed(-14, 8),
    to_signed(-13, 8),
    to_signed(-10, 8),
    to_signed(-4, 8),
    to_signed(1, 8),
    to_signed(4, 8),
    to_signed(6, 8),
    to_signed(5, 8),
    to_signed(1, 8),
    to_signed(-5, 8),
    to_signed(-11, 8),
    to_signed(-15, 8),
    to_signed(-17, 8),
    to_signed(-18, 8),
    to_signed(-16, 8),
    to_signed(-10, 8),
    to_signed(1, 8),
    to_signed(16, 8),
    to_signed(33, 8),
    to_signed(49, 8),
    to_signed(59, 8),
    to_signed(61, 8),
    to_signed(57, 8),
    to_signed(51, 8),
    to_signed(43, 8),
    to_signed(34, 8),
    to_signed(27, 8),
    to_signed(21, 8),
    to_signed(16, 8),
    to_signed(13, 8),
    to_signed(14, 8),
    to_signed(17, 8),
    to_signed(21, 8),
    to_signed(25, 8),
    to_signed(29, 8),
    to_signed(33, 8),
    to_signed(36, 8),
    to_signed(40, 8),
    to_signed(41, 8),
    to_signed(38, 8),
    to_signed(29, 8),
    to_signed(18, 8),
    to_signed(1, 8),
    to_signed(-20, 8),
    to_signed(-44, 8),
    to_signed(-65, 8),
    to_signed(-80, 8),
    to_signed(-85, 8),
    to_signed(-77, 8),
    to_signed(-57, 8),
    to_signed(-31, 8),
    to_signed(-5, 8),
    to_signed(15, 8),
    to_signed(28, 8),
    to_signed(29, 8),
    to_signed(17, 8),
    to_signed(-3, 8),
    to_signed(-23, 8),
    to_signed(-38, 8),
    to_signed(-49, 8),
    to_signed(-52, 8),
    to_signed(-45, 8),
    to_signed(-29, 8),
    to_signed(-10, 8),
    to_signed(9, 8),
    to_signed(24, 8),
    to_signed(32, 8),
    to_signed(32, 8),
    to_signed(27, 8),
    to_signed(18, 8),
    to_signed(7, 8),
    to_signed(-5, 8),
    to_signed(-13, 8),
    to_signed(-16, 8),
    to_signed(-16, 8),
    to_signed(-13, 8),
    to_signed(-7, 8),
    to_signed(1, 8),
    to_signed(6, 8),
    to_signed(8, 8),
    to_signed(9, 8),
    to_signed(9, 8),
    to_signed(5, 8),
    to_signed(0, 8),
    to_signed(-4, 8),
    to_signed(-7, 8),
    to_signed(-9, 8),
    to_signed(-8, 8),
    to_signed(-3, 8),
    to_signed(4, 8),
    to_signed(14, 8),
    to_signed(27, 8),
    to_signed(40, 8),
    to_signed(46, 8),
    to_signed(45, 8),
    to_signed(39, 8),
    to_signed(32, 8),
    to_signed(24, 8),
    to_signed(15, 8),
    to_signed(6, 8),
    to_signed(0, 8),
    to_signed(-2, 8),
    to_signed(-1, 8),
    to_signed(4, 8),
    to_signed(11, 8),
    to_signed(17, 8),
    to_signed(21, 8),
    to_signed(26, 8),
    to_signed(33, 8),
    to_signed(37, 8),
    to_signed(38, 8),
    to_signed(36, 8),
    to_signed(34, 8),
    to_signed(28, 8),
    to_signed(15, 8),
    to_signed(-3, 8),
    to_signed(-22, 8),
    to_signed(-43, 8),
    to_signed(-67, 8),
    to_signed(-86, 8),
    to_signed(-93, 8),
    to_signed(-87, 8),
    to_signed(-71, 8),
    to_signed(-47, 8),
    to_signed(-21, 8),
    to_signed(1, 8),
    to_signed(15, 8),
    to_signed(19, 8),
    to_signed(13, 8),
    to_signed(-2, 8),
    to_signed(-20, 8),
    to_signed(-38, 8),
    to_signed(-51, 8),
    to_signed(-59, 8),
    to_signed(-58, 8),
    to_signed(-47, 8),
    to_signed(-30, 8),
    to_signed(-10, 8),
    to_signed(10, 8),
    to_signed(24, 8),
    to_signed(29, 8),
    to_signed(27, 8),
    to_signed(20, 8),
    to_signed(12, 8),
    to_signed(1, 8),
    to_signed(-11, 8),
    to_signed(-19, 8),
    to_signed(-23, 8),
    to_signed(-23, 8),
    to_signed(-19, 8),
    to_signed(-12, 8),
    to_signed(-6, 8),
    to_signed(-2, 8),
    to_signed(0, 8),
    to_signed(-1, 8),
    to_signed(-5, 8),
    to_signed(-12, 8),
    to_signed(-20, 8),
    to_signed(-27, 8),
    to_signed(-31, 8),
    to_signed(-28, 8),
    to_signed(-20, 8),
    to_signed(-7, 8),
    to_signed(8, 8),
    to_signed(20, 8),
    to_signed(28, 8),
    to_signed(33, 8),
    to_signed(33, 8),
    to_signed(30, 8),
    to_signed(24, 8),
    to_signed(16, 8),
    to_signed(8, 8),
    to_signed(1, 8),
    to_signed(-3, 8),
    to_signed(-2, 8),
    to_signed(1, 8),
    to_signed(6, 8),
    to_signed(10, 8),
    to_signed(14, 8),
    to_signed(18, 8),
    to_signed(22, 8),
    to_signed(27, 8),
    to_signed(32, 8),
    to_signed(34, 8),
    to_signed(33, 8),
    to_signed(29, 8),
    to_signed(21, 8),
    to_signed(7, 8),
    to_signed(-11, 8),
    to_signed(-30, 8),
    to_signed(-51, 8),
    to_signed(-71, 8),
    to_signed(-84, 8),
    to_signed(-86, 8),
    to_signed(-77, 8),
    to_signed(-59, 8),
    to_signed(-35, 8),
    to_signed(-10, 8),
    to_signed(11, 8),
    to_signed(23, 8),
    to_signed(24, 8),
    to_signed(16, 8),
    to_signed(-2, 8),
    to_signed(-24, 8),
    to_signed(-45, 8),
    to_signed(-60, 8),
    to_signed(-68, 8),
    to_signed(-65, 8),
    to_signed(-51, 8),
    to_signed(-29, 8),
    to_signed(-7, 8),
    to_signed(12, 8),
    to_signed(26, 8),
    to_signed(33, 8),
    to_signed(30, 8),
    to_signed(19, 8),
    to_signed(6, 8),
    to_signed(-6, 8),
    to_signed(-17, 8),
    to_signed(-22, 8),
    to_signed(-20, 8),
    to_signed(-17, 8),
    to_signed(-13, 8),
    to_signed(-7, 8),
    to_signed(1, 8),
    to_signed(7, 8),
    to_signed(8, 8),
    to_signed(6, 8),
    to_signed(2, 8),
    to_signed(-2, 8),
    to_signed(-7, 8),
    to_signed(-12, 8),
    to_signed(-13, 8),
    to_signed(-10, 8),
    to_signed(-3, 8),
    to_signed(8, 8),
    to_signed(21, 8),
    to_signed(31, 8),
    to_signed(39, 8),
    to_signed(47, 8),
    to_signed(56, 8),
    to_signed(59, 8),
    to_signed(57, 8),
    to_signed(51, 8),
    to_signed(42, 8),
    to_signed(30, 8),
    to_signed(17, 8),
    to_signed(7, 8),
    to_signed(4, 8),
    to_signed(7, 8),
    to_signed(16, 8),
    to_signed(28, 8),
    to_signed(40, 8),
    to_signed(50, 8),
    to_signed(58, 8),
    to_signed(61, 8),
    to_signed(59, 8),
    to_signed(52, 8),
    to_signed(41, 8),
    to_signed(28, 8),
    to_signed(12, 8),
    to_signed(-6, 8),
    to_signed(-24, 8),
    to_signed(-42, 8),
    to_signed(-55, 8),
    to_signed(-63, 8),
    to_signed(-62, 8),
    to_signed(-50, 8),
    to_signed(-30, 8),
    to_signed(-7, 8),
    to_signed(12, 8),
    to_signed(25, 8),
    to_signed(28, 8),
    to_signed(20, 8),
    to_signed(4, 8),
    to_signed(-16, 8),
    to_signed(-36, 8),
    to_signed(-54, 8),
    to_signed(-65, 8),
    to_signed(-65, 8),
    to_signed(-55, 8),
    to_signed(-37, 8),
    to_signed(-16, 8),
    to_signed(5, 8),
    to_signed(19, 8),
    to_signed(27, 8),
    to_signed(30, 8),
    to_signed(25, 8),
    to_signed(14, 8),
    to_signed(0, 8),
    to_signed(-10, 8),
    to_signed(-18, 8),
    to_signed(-25, 8),
    to_signed(-28, 8),
    to_signed(-25, 8),
    to_signed(-18, 8),
    to_signed(-9, 8),
    to_signed(0, 8),
    to_signed(9, 8),
    to_signed(16, 8),
    to_signed(17, 8),
    to_signed(12, 8),
    to_signed(3, 8),
    to_signed(-7, 8),
    to_signed(-12, 8),
    to_signed(-11, 8),
    to_signed(-6, 8),
    to_signed(3, 8),
    to_signed(16, 8),
    to_signed(30, 8),
    to_signed(39, 8),
    to_signed(44, 8),
    to_signed(46, 8),
    to_signed(45, 8),
    to_signed(42, 8),
    to_signed(36, 8),
    to_signed(29, 8),
    to_signed(20, 8),
    to_signed(11, 8),
    to_signed(1, 8),
    to_signed(-6, 8),
    to_signed(-7, 8),
    to_signed(-2, 8),
    to_signed(10, 8),
    to_signed(26, 8),
    to_signed(41, 8),
    to_signed(52, 8),
    to_signed(56, 8),
    to_signed(56, 8),
    to_signed(51, 8),
    to_signed(42, 8),
    to_signed(30, 8),
    to_signed(16, 8),
    to_signed(2, 8),
    to_signed(-11, 8),
    to_signed(-25, 8),
    to_signed(-40, 8),
    to_signed(-54, 8),
    to_signed(-64, 8),
    to_signed(-68, 8),
    to_signed(-63, 8),
    to_signed(-48, 8),
    to_signed(-27, 8),
    to_signed(-4, 8),
    to_signed(17, 8),
    to_signed(27, 8),
    to_signed(24, 8),
    to_signed(8, 8),
    to_signed(-13, 8),
    to_signed(-37, 8),
    to_signed(-60, 8),
    to_signed(-77, 8),
    to_signed(-81, 8),
    to_signed(-72, 8),
    to_signed(-52, 8),
    to_signed(-26, 8),
    to_signed(1, 8),
    to_signed(21, 8),
    to_signed(28, 8),
    to_signed(27, 8),
    to_signed(20, 8),
    to_signed(10, 8),
    to_signed(-2, 8),
    to_signed(-13, 8),
    to_signed(-21, 8),
    to_signed(-24, 8),
    to_signed(-22, 8),
    to_signed(-17, 8),
    to_signed(-12, 8),
    to_signed(-8, 8),
    to_signed(-5, 8),
    to_signed(0, 8),
    to_signed(4, 8),
    to_signed(3, 8),
    to_signed(-1, 8),
    to_signed(-4, 8),
    to_signed(-4, 8),
    to_signed(-5, 8),
    to_signed(-7, 8),
    to_signed(-5, 8),
    to_signed(1, 8),
    to_signed(10, 8),
    to_signed(19, 8),
    to_signed(26, 8),
    to_signed(31, 8),
    to_signed(33, 8),
    to_signed(35, 8),
    to_signed(35, 8),
    to_signed(33, 8),
    to_signed(28, 8),
    to_signed(21, 8),
    to_signed(13, 8),
    to_signed(6, 8),
    to_signed(5, 8),
    to_signed(9, 8),
    to_signed(17, 8),
    to_signed(26, 8),
    to_signed(33, 8),
    to_signed(41, 8),
    to_signed(49, 8),
    to_signed(54, 8),
    to_signed(52, 8),
    to_signed(44, 8),
    to_signed(33, 8),
    to_signed(21, 8),
    to_signed(8, 8),
    to_signed(-6, 8),
    to_signed(-22, 8),
    to_signed(-40, 8),
    to_signed(-57, 8),
    to_signed(-69, 8),
    to_signed(-71, 8),
    to_signed(-63, 8),
    to_signed(-45, 8),
    to_signed(-20, 8),
    to_signed(5, 8),
    to_signed(21, 8),
    to_signed(26, 8),
    to_signed(20, 8),
    to_signed(5, 8),
    to_signed(-16, 8),
    to_signed(-39, 8),
    to_signed(-57, 8),
    to_signed(-66, 8),
    to_signed(-63, 8),
    to_signed(-51, 8),
    to_signed(-33, 8),
    to_signed(-10, 8),
    to_signed(10, 8),
    to_signed(24, 8),
    to_signed(29, 8),
    to_signed(26, 8),
    to_signed(18, 8),
    to_signed(7, 8),
    to_signed(-3, 8),
    to_signed(-9, 8),
    to_signed(-13, 8),
    to_signed(-14, 8),
    to_signed(-13, 8),
    to_signed(-14, 8),
    to_signed(-14, 8),
    to_signed(-11, 8),
    to_signed(-5, 8),
    to_signed(2, 8),
    to_signed(6, 8),
    to_signed(8, 8),
    to_signed(7, 8),
    to_signed(0, 8),
    to_signed(-9, 8),
    to_signed(-17, 8),
    to_signed(-22, 8),
    to_signed(-20, 8),
    to_signed(-13, 8),
    to_signed(-2, 8),
    to_signed(10, 8),
    to_signed(22, 8),
    to_signed(33, 8),
    to_signed(42, 8),
    to_signed(46, 8),
    to_signed(45, 8),
    to_signed(40, 8),
    to_signed(33, 8),
    to_signed(22, 8),
    to_signed(10, 8),
    to_signed(-1, 8),
    to_signed(-6, 8),
    to_signed(-5, 8),
    to_signed(1, 8),
    to_signed(10, 8),
    to_signed(20, 8),
    to_signed(30, 8),
    to_signed(40, 8),
    to_signed(47, 8),
    to_signed(52, 8),
    to_signed(52, 8),
    to_signed(46, 8),
    to_signed(34, 8),
    to_signed(17, 8),
    to_signed(-3, 8),
    to_signed(-23, 8),
    to_signed(-41, 8),
    to_signed(-56, 8),
    to_signed(-67, 8),
    to_signed(-70, 8),
    to_signed(-65, 8),
    to_signed(-51, 8),
    to_signed(-33, 8),
    to_signed(-12, 8),
    to_signed(6, 8),
    to_signed(18, 8),
    to_signed(19, 8),
    to_signed(12, 8),
    to_signed(-2, 8),
    to_signed(-21, 8),
    to_signed(-42, 8),
    to_signed(-60, 8),
    to_signed(-71, 8),
    to_signed(-71, 8),
    to_signed(-60, 8),
    to_signed(-40, 8),
    to_signed(-16, 8),
    to_signed(5, 8),
    to_signed(20, 8),
    to_signed(28, 8),
    to_signed(29, 8),
    to_signed(21, 8),
    to_signed(8, 8),
    to_signed(-4, 8),
    to_signed(-12, 8),
    to_signed(-17, 8),
    to_signed(-21, 8),
    to_signed(-22, 8),
    to_signed(-19, 8),
    to_signed(-14, 8),
    to_signed(-8, 8),
    to_signed(0, 8),
    to_signed(7, 8),
    to_signed(10, 8),
    to_signed(11, 8),
    to_signed(7, 8),
    to_signed(-1, 8),
    to_signed(-10, 8),
    to_signed(-16, 8),
    to_signed(-16, 8),
    to_signed(-10, 8),
    to_signed(0, 8),
    to_signed(13, 8),
    to_signed(26, 8),
    to_signed(38, 8),
    to_signed(44, 8),
    to_signed(46, 8),
    to_signed(45, 8),
    to_signed(41, 8),
    to_signed(35, 8),
    to_signed(27, 8),
    to_signed(20, 8),
    to_signed(16, 8),
    to_signed(16, 8),
    to_signed(16, 8),
    to_signed(17, 8),
    to_signed(18, 8),
    to_signed(20, 8),
    to_signed(25, 8),
    to_signed(31, 8),
    to_signed(38, 8),
    to_signed(44, 8),
    to_signed(51, 8),
    to_signed(57, 8),
    to_signed(56, 8),
    to_signed(46, 8),
    to_signed(32, 8),
    to_signed(16, 8),
    to_signed(-2, 8),
    to_signed(-25, 8),
    to_signed(-49, 8),
    to_signed(-68, 8),
    to_signed(-75, 8),
    to_signed(-69, 8),
    to_signed(-55, 8),
    to_signed(-36, 8),
    to_signed(-15, 8),
    to_signed(4, 8),
    to_signed(18, 8),
    to_signed(23, 8),
    to_signed(16, 8),
    to_signed(0, 8),
    to_signed(-19, 8),
    to_signed(-40, 8),
    to_signed(-59, 8),
    to_signed(-71, 8),
    to_signed(-72, 8),
    to_signed(-64, 8),
    to_signed(-48, 8),
    to_signed(-27, 8),
    to_signed(-6, 8),
    to_signed(9, 8),
    to_signed(18, 8),
    to_signed(21, 8),
    to_signed(18, 8),
    to_signed(10, 8),
    to_signed(-1, 8),
    to_signed(-11, 8),
    to_signed(-18, 8),
    to_signed(-23, 8),
    to_signed(-25, 8),
    to_signed(-24, 8),
    to_signed(-20, 8),
    to_signed(-13, 8),
    to_signed(-2, 8),
    to_signed(7, 8),
    to_signed(13, 8),
    to_signed(15, 8),
    to_signed(13, 8),
    to_signed(8, 8),
    to_signed(1, 8),
    to_signed(-6, 8),
    to_signed(-9, 8),
    to_signed(-8, 8),
    to_signed(-5, 8),
    to_signed(0, 8),
    to_signed(5, 8),
    to_signed(11, 8),
    to_signed(14, 8),
    to_signed(15, 8),
    to_signed(18, 8),
    to_signed(22, 8),
    to_signed(24, 8),
    to_signed(22, 8),
    to_signed(16, 8),
    to_signed(9, 8),
    to_signed(4, 8),
    to_signed(0, 8),
    to_signed(-2, 8),
    to_signed(-3, 8),
    to_signed(1, 8),
    to_signed(8, 8),
    to_signed(17, 8),
    to_signed(25, 8),
    to_signed(32, 8),
    to_signed(39, 8),
    to_signed(45, 8),
    to_signed(46, 8),
    to_signed(41, 8),
    to_signed(32, 8),
    to_signed(19, 8),
    to_signed(1, 8),
    to_signed(-20, 8),
    to_signed(-39, 8),
    to_signed(-55, 8),
    to_signed(-66, 8),
    to_signed(-71, 8),
    to_signed(-66, 8),
    to_signed(-50, 8),
    to_signed(-28, 8),
    to_signed(-7, 8),
    to_signed(10, 8),
    to_signed(22, 8),
    to_signed(25, 8),
    to_signed(17, 8),
    to_signed(-1, 8),
    to_signed(-23, 8),
    to_signed(-44, 8),
    to_signed(-60, 8),
    to_signed(-69, 8),
    to_signed(-71, 8),
    to_signed(-63, 8),
    to_signed(-47, 8),
    to_signed(-25, 8),
    to_signed(-5, 8),
    to_signed(9, 8),
    to_signed(16, 8),
    to_signed(18, 8),
    to_signed(14, 8),
    to_signed(4, 8),
    to_signed(-7, 8),
    to_signed(-16, 8),
    to_signed(-22, 8),
    to_signed(-25, 8),
    to_signed(-25, 8),
    to_signed(-21, 8),
    to_signed(-15, 8),
    to_signed(-8, 8),
    to_signed(0, 8),
    to_signed(9, 8),
    to_signed(16, 8),
    to_signed(20, 8),
    to_signed(20, 8),
    to_signed(15, 8),
    to_signed(6, 8),
    to_signed(-4, 8),
    to_signed(-8, 8),
    to_signed(-6, 8),
    to_signed(-2, 8),
    to_signed(5, 8),
    to_signed(13, 8),
    to_signed(22, 8),
    to_signed(30, 8),
    to_signed(37, 8),
    to_signed(45, 8),
    to_signed(51, 8),
    to_signed(54, 8),
    to_signed(54, 8),
    to_signed(52, 8),
    to_signed(45, 8),
    to_signed(37, 8),
    to_signed(30, 8),
    to_signed(28, 8),
    to_signed(26, 8),
    to_signed(26, 8),
    to_signed(30, 8),
    to_signed(37, 8),
    to_signed(45, 8),
    to_signed(51, 8),
    to_signed(54, 8),
    to_signed(55, 8),
    to_signed(53, 8),
    to_signed(48, 8),
    to_signed(41, 8),
    to_signed(29, 8),
    to_signed(13, 8),
    to_signed(-5, 8),
    to_signed(-23, 8),
    to_signed(-37, 8),
    to_signed(-45, 8),
    to_signed(-44, 8),
    to_signed(-32, 8),
    to_signed(-13, 8),
    to_signed(5, 8),
    to_signed(20, 8),
    to_signed(29, 8),
    to_signed(31, 8),
    to_signed(22, 8),
    to_signed(6, 8),
    to_signed(-14, 8),
    to_signed(-33, 8),
    to_signed(-47, 8),
    to_signed(-56, 8),
    to_signed(-56, 8),
    to_signed(-47, 8),
    to_signed(-31, 8),
    to_signed(-11, 8),
    to_signed(6, 8),
    to_signed(16, 8),
    to_signed(19, 8),
    to_signed(19, 8),
    to_signed(15, 8),
    to_signed(7, 8),
    to_signed(-2, 8),
    to_signed(-9, 8),
    to_signed(-12, 8),
    to_signed(-16, 8),
    to_signed(-22, 8),
    to_signed(-25, 8),
    to_signed(-24, 8),
    to_signed(-19, 8),
    to_signed(-13, 8),
    to_signed(-4, 8),
    to_signed(8, 8),
    to_signed(18, 8),
    to_signed(21, 8),
    to_signed(19, 8),
    to_signed(12, 8),
    to_signed(4, 8),
    to_signed(-3, 8),
    to_signed(-6, 8),
    to_signed(-5, 8),
    to_signed(-1, 8),
    to_signed(4, 8),
    to_signed(10, 8),
    to_signed(16, 8),
    to_signed(22, 8),
    to_signed(28, 8),
    to_signed(34, 8),
    to_signed(36, 8),
    to_signed(34, 8),
    to_signed(31, 8),
    to_signed(27, 8),
    to_signed(21, 8),
    to_signed(14, 8),
    to_signed(9, 8),
    to_signed(7, 8),
    to_signed(7, 8),
    to_signed(10, 8),
    to_signed(15, 8),
    to_signed(21, 8),
    to_signed(27, 8),
    to_signed(32, 8),
    to_signed(35, 8),
    to_signed(35, 8),
    to_signed(29, 8),
    to_signed(18, 8),
    to_signed(5, 8),
    to_signed(-6, 8),
    to_signed(-16, 8),
    to_signed(-26, 8),
    to_signed(-33, 8),
    to_signed(-36, 8),
    to_signed(-35, 8),
    to_signed(-29, 8),
    to_signed(-21, 8),
    to_signed(-11, 8),
    to_signed(-3, 8),
    to_signed(3, 8),
    to_signed(5, 8),
    to_signed(1, 8),
    to_signed(-7, 8),
    to_signed(-17, 8),
    to_signed(-29, 8),
    to_signed(-40, 8),
    to_signed(-48, 8),
    to_signed(-49, 8),
    to_signed(-45, 8),
    to_signed(-38, 8),
    to_signed(-28, 8),
    to_signed(-17, 8),
    to_signed(-5, 8),
    to_signed(4, 8),
    to_signed(6, 8),
    to_signed(1, 8),
    to_signed(-7, 8),
    to_signed(-15, 8),
    to_signed(-22, 8),
    to_signed(-27, 8),
    to_signed(-29, 8),
    to_signed(-30, 8),
    to_signed(-30, 8),
    to_signed(-30, 8),
    to_signed(-26, 8),
    to_signed(-19, 8),
    to_signed(-8, 8),
    to_signed(2, 8),
    to_signed(6, 8),
    to_signed(5, 8),
    to_signed(2, 8),
    to_signed(-1, 8),
    to_signed(-5, 8),
    to_signed(-9, 8),
    to_signed(-10, 8),
    to_signed(-8, 8),
    to_signed(-5, 8),
    to_signed(-4, 8),
    to_signed(-4, 8),
    to_signed(-4, 8),
    to_signed(-2, 8),
    to_signed(2, 8),
    to_signed(6, 8),
    to_signed(8, 8),
    to_signed(9, 8),
    to_signed(10, 8),
    to_signed(11, 8),
    to_signed(10, 8),
    to_signed(6, 8),
    to_signed(2, 8),
    to_signed(1, 8),
    to_signed(2, 8),
    to_signed(4, 8),
    to_signed(4, 8),
    to_signed(7, 8),
    to_signed(12, 8),
    to_signed(16, 8),
    to_signed(18, 8),
    to_signed(16, 8),
    to_signed(13, 8),
    to_signed(9, 8),
    to_signed(4, 8),
    to_signed(-1, 8),
    to_signed(-4, 8),
    to_signed(-5, 8),
    to_signed(-5, 8),
    to_signed(-6, 8),
    to_signed(-10, 8),
    to_signed(-13, 8),
    to_signed(-15, 8),
    to_signed(-13, 8),
    to_signed(-10, 8),
    to_signed(-6, 8),
    to_signed(-1, 8),
    to_signed(2, 8),
    to_signed(3, 8),
    to_signed(-1, 8),
    to_signed(-5, 8),
    to_signed(-10, 8),
    to_signed(-13, 8),
    to_signed(-14, 8),
    to_signed(-12, 8),
    to_signed(-8, 8),
    to_signed(-4, 8),
    to_signed(0, 8),
    to_signed(3, 8),
    to_signed(6, 8),
    to_signed(9, 8),
    to_signed(10, 8),
    to_signed(9, 8),
    to_signed(7, 8),
    to_signed(4, 8),
    to_signed(2, 8),
    to_signed(3, 8),
    to_signed(4, 8),
    to_signed(4, 8),
    to_signed(4, 8),
    to_signed(5, 8),
    to_signed(6, 8),
    to_signed(6, 8),
    to_signed(6, 8),
    to_signed(6, 8),
    to_signed(7, 8),
    to_signed(9, 8),
    to_signed(9, 8),
    to_signed(8, 8),
    to_signed(6, 8),
    to_signed(5, 8),
    to_signed(2, 8),
    to_signed(-2, 8),
    to_signed(-7, 8),
    to_signed(-9, 8),
    to_signed(-11, 8),
    to_signed(-11, 8),
    to_signed(-9, 8),
    to_signed(-5, 8),
    to_signed(2, 8),
    to_signed(8, 8),
    to_signed(12, 8),
    to_signed(13, 8),
    to_signed(11, 8),
    to_signed(8, 8),
    to_signed(5, 8),
    to_signed(3, 8),
    to_signed(1, 8),
    to_signed(0, 8),
    to_signed(3, 8),
    to_signed(5, 8),
    to_signed(6, 8),
    to_signed(6, 8),
    to_signed(6, 8),
    to_signed(6, 8),
    to_signed(5, 8),
    to_signed(2, 8),
    to_signed(0, 8),
    to_signed(-1, 8),
    to_signed(-3, 8),
    to_signed(-6, 8),
    to_signed(-10, 8),
    to_signed(-12, 8),
    to_signed(-12, 8),
    to_signed(-13, 8),
    to_signed(-13, 8),
    to_signed(-11, 8),
    to_signed(-7, 8),
    to_signed(-2, 8),
    to_signed(0, 8),
    to_signed(-2, 8),
    to_signed(-8, 8),
    to_signed(-14, 8),
    to_signed(-19, 8),
    to_signed(-21, 8),
    to_signed(-20, 8),
    to_signed(-16, 8),
    to_signed(-11, 8),
    to_signed(-6, 8),
    to_signed(-2, 8),
    to_signed(-1, 8),
    to_signed(1, 8),
    to_signed(3, 8),
    to_signed(6, 8),
    to_signed(6, 8),
    to_signed(3, 8),
    to_signed(-2, 8),
    to_signed(-5, 8),
    to_signed(-5, 8),
    to_signed(-3, 8),
    to_signed(-1, 8),
    to_signed(0, 8),
    to_signed(0, 8),
    to_signed(2, 8),
    to_signed(2, 8),
    to_signed(-1, 8),
    to_signed(-4, 8),
    to_signed(-3, 8),
    to_signed(1, 8),
    to_signed(4, 8),
    to_signed(6, 8),
    to_signed(7, 8),
    to_signed(8, 8),
    to_signed(7, 8),
    to_signed(3, 8),
    to_signed(-2, 8),
    to_signed(-6, 8),
    to_signed(-10, 8),
    to_signed(-13, 8),
    to_signed(-14, 8),
    to_signed(-12, 8),
    to_signed(-8, 8),
    to_signed(-2, 8),
    to_signed(4, 8),
    to_signed(9, 8),
    to_signed(11, 8),
    to_signed(9, 8),
    to_signed(6, 8),
    to_signed(3, 8),
    to_signed(2, 8),
    to_signed(1, 8),
    to_signed(3, 8),
    to_signed(6, 8),
    to_signed(8, 8),
    to_signed(10, 8),
    to_signed(11, 8),
    to_signed(11, 8),
    to_signed(9, 8),
    to_signed(8, 8),
    to_signed(7, 8),
    to_signed(6, 8),
    to_signed(2, 8),
    to_signed(-1, 8),
    to_signed(-3, 8),
    to_signed(-3, 8),
    to_signed(-4, 8),
    to_signed(-7, 8),
    to_signed(-8, 8),
    to_signed(-7, 8),
    to_signed(-6, 8),
    to_signed(-6, 8),
    to_signed(-7, 8),
    to_signed(-7, 8),
    to_signed(-6, 8),
    to_signed(-6, 8),
    to_signed(-7, 8),
    to_signed(-8, 8),
    to_signed(-5, 8),
    to_signed(-2, 8),
    to_signed(-4, 8),
    to_signed(-10, 8),
    to_signed(-13, 8),
    to_signed(-10, 8),
    to_signed(-3, 8),
    to_signed(1, 8),
    to_signed(1, 8),
    to_signed(3, 8),
    to_signed(7, 8),
    to_signed(10, 8),
    to_signed(8, 8),
    to_signed(4, 8),
    to_signed(0, 8),
    to_signed(-1, 8),
    to_signed(0, 8),
    to_signed(1, 8),
    to_signed(3, 8),
    to_signed(6, 8),
    to_signed(9, 8),
    to_signed(12, 8),
    to_signed(14, 8),
    to_signed(16, 8),
    to_signed(17, 8),
    to_signed(17, 8),
    to_signed(17, 8),
    to_signed(18, 8),
    to_signed(17, 8),
    to_signed(15, 8),
    to_signed(11, 8),
    to_signed(7, 8),
    to_signed(4, 8),
    to_signed(2, 8),
    to_signed(0, 8),
    to_signed(-3, 8),
    to_signed(-5, 8),
    to_signed(-7, 8),
    to_signed(-5, 8),
    to_signed(-2, 8),
    to_signed(2, 8),
    to_signed(4, 8),
    to_signed(5, 8),
    to_signed(4, 8),
    to_signed(3, 8),
    to_signed(1, 8),
    to_signed(-1, 8),
    to_signed(-1, 8),
    to_signed(0, 8),
    to_signed(0, 8),
    to_signed(1, 8),
    to_signed(2, 8),
    to_signed(3, 8),
    to_signed(2, 8),
    to_signed(2, 8),
    to_signed(3, 8),
    to_signed(2, 8),
    to_signed(-2, 8),
    to_signed(-6, 8),
    to_signed(-8, 8),
    to_signed(-8, 8),
    to_signed(-7, 8),
    to_signed(-5, 8),
    to_signed(-3, 8),
    to_signed(-2, 8),
    to_signed(-2, 8),
    to_signed(-1, 8),
    to_signed(-2, 8),
    to_signed(-3, 8),
    to_signed(-5, 8),
    to_signed(-8, 8),
    to_signed(-9, 8),
    to_signed(-10, 8),
    to_signed(-9, 8),
    to_signed(-7, 8),
    to_signed(-5, 8),
    to_signed(-5, 8),
    to_signed(-5, 8),
    to_signed(-4, 8),
    to_signed(-4, 8),
    to_signed(-5, 8),
    to_signed(-5, 8),
    to_signed(-5, 8),
    to_signed(-3, 8),
    to_signed(-1, 8),
    to_signed(0, 8),
    to_signed(0, 8),
    to_signed(1, 8),
    to_signed(4, 8),
    to_signed(6, 8),
    to_signed(5, 8),
    to_signed(2, 8),
    to_signed(3, 8),
    to_signed(7, 8),
    to_signed(11, 8),
    to_signed(13, 8),
    to_signed(13, 8),
    to_signed(14, 8),
    to_signed(14, 8),
    to_signed(14, 8),
    to_signed(11, 8),
    to_signed(7, 8),
    to_signed(5, 8),
    to_signed(4, 8),
    to_signed(3, 8),
    to_signed(-1, 8),
    to_signed(-6, 8),
    to_signed(-9, 8),
    to_signed(-12, 8),
    to_signed(-13, 8),
    to_signed(-11, 8),
    to_signed(-5, 8),
    to_signed(0, 8),
    to_signed(4, 8),
    to_signed(5, 8),
    to_signed(5, 8),
    to_signed(3, 8),
    to_signed(1, 8),
    to_signed(0, 8),
    to_signed(0, 8),
    to_signed(0, 8),
    to_signed(0, 8),
    to_signed(-1, 8),
    to_signed(0, 8),
    to_signed(2, 8),
    to_signed(1, 8),
    to_signed(-2, 8),
    to_signed(-4, 8),
    to_signed(-6, 8),
    to_signed(-7, 8),
    to_signed(-8, 8),
    to_signed(-8, 8),
    to_signed(-7, 8),
    to_signed(-6, 8),
    to_signed(-4, 8),
    to_signed(-2, 8),
    to_signed(-2, 8),
    to_signed(-2, 8),
    to_signed(-2, 8),
    to_signed(-2, 8),
    to_signed(-3, 8),
    to_signed(-4, 8),
    to_signed(-6, 8),
    to_signed(-8, 8),
    to_signed(-9, 8),
    to_signed(-10, 8),
    to_signed(-11, 8),
    to_signed(-13, 8),
    to_signed(-13, 8),
    to_signed(-12, 8),
    to_signed(-9, 8),
    to_signed(-4, 8),
    to_signed(-1, 8),
    to_signed(0, 8),
    to_signed(-1, 8),
    to_signed(0, 8),
    to_signed(2, 8),
    to_signed(5, 8),
    to_signed(8, 8),
    to_signed(8, 8),
    to_signed(6, 8),
    to_signed(2, 8),
    to_signed(-1, 8),
    to_signed(-3, 8),
    to_signed(-3, 8),
    to_signed(-1, 8),
    to_signed(1, 8),
    to_signed(1, 8),
    to_signed(-1, 8),
    to_signed(-1, 8),
    to_signed(0, 8),
    to_signed(0, 8),
    to_signed(-1, 8),
    to_signed(0, 8),
    to_signed(1, 8),
    to_signed(2, 8),
    to_signed(1, 8),
    to_signed(-2, 8),
    to_signed(-5, 8),
    to_signed(-10, 8),
    to_signed(-14, 8),
    to_signed(-18, 8),
    to_signed(-20, 8),
    to_signed(-19, 8),
    to_signed(-17, 8),
    to_signed(-14, 8),
    to_signed(-12, 8),
    to_signed(-9, 8),
    to_signed(-7, 8),
    to_signed(-3, 8),
    to_signed(1, 8),
    to_signed(3, 8),
    to_signed(2, 8),
    to_signed(-1, 8),
    to_signed(-3, 8),
    to_signed(-4, 8),
    to_signed(-4, 8),
    to_signed(-3, 8),
    to_signed(-2, 8),
    to_signed(0, 8),
    to_signed(1, 8),
    to_signed(-2, 8),
    to_signed(-7, 8),
    to_signed(-12, 8),
    to_signed(-14, 8),
    to_signed(-15, 8),
    to_signed(-15, 8),
    to_signed(-13, 8),
    to_signed(-11, 8),
    to_signed(-9, 8),
    to_signed(-9, 8),
    to_signed(-9, 8),
    to_signed(-7, 8),
    to_signed(-6, 8),
    to_signed(-7, 8),
    to_signed(-10, 8),
    to_signed(-13, 8),
    to_signed(-15, 8),
    to_signed(-15, 8),
    to_signed(-15, 8),
    to_signed(-15, 8),
    to_signed(-14, 8),
    to_signed(-13, 8),
    to_signed(-13, 8),
    to_signed(-15, 8),
    to_signed(-17, 8),
    to_signed(-16, 8),
    to_signed(-12, 8),
    to_signed(-8, 8),
    to_signed(-5, 8),
    to_signed(-3, 8),
    to_signed(-2, 8),
    to_signed(-3, 8),
    to_signed(-4, 8),
    to_signed(-6, 8),
    to_signed(-6, 8),
    to_signed(-3, 8),
    to_signed(-1, 8),
    to_signed(-2, 8),
    to_signed(-3, 8),
    to_signed(-3, 8),
    to_signed(-1, 8),
    to_signed(-1, 8),
    to_signed(-2, 8),
    to_signed(-3, 8),
    to_signed(-2, 8),
    to_signed(0, 8),
    to_signed(1, 8),
    to_signed(0, 8),
    to_signed(1, 8),
    to_signed(2, 8),
    to_signed(4, 8),
    to_signed(4, 8),
    to_signed(4, 8),
    to_signed(1, 8),
    to_signed(-1, 8),
    to_signed(-2, 8),
    to_signed(-1, 8),
    to_signed(1, 8),
    to_signed(5, 8),
    to_signed(8, 8),
    to_signed(9, 8),
    to_signed(11, 8),
    to_signed(14, 8),
    to_signed(14, 8),
    to_signed(11, 8),
    to_signed(9, 8),
    to_signed(9, 8),
    to_signed(9, 8),
    to_signed(7, 8),
    to_signed(5, 8),
    to_signed(7, 8),
    to_signed(12, 8),
    to_signed(14, 8),
    to_signed(13, 8),
    to_signed(10, 8),
    to_signed(7, 8),
    to_signed(3, 8),
    to_signed(-1, 8),
    to_signed(-4, 8),
    to_signed(-4, 8),
    to_signed(0, 8),
    to_signed(4, 8),
    to_signed(7, 8),
    to_signed(8, 8),
    to_signed(7, 8),
    to_signed(5, 8),
    to_signed(2, 8),
    to_signed(-1, 8),
    to_signed(-3, 8),
    to_signed(-2, 8),
    to_signed(0, 8),
    to_signed(1, 8),
    to_signed(2, 8),
    to_signed(2, 8),
    to_signed(4, 8),
    to_signed(7, 8),
    to_signed(8, 8),
    to_signed(8, 8),
    to_signed(6, 8),
    to_signed(5, 8),
    to_signed(6, 8),
    to_signed(8, 8),
    to_signed(8, 8),
    to_signed(10, 8),
    to_signed(11, 8),
    to_signed(12, 8),
    to_signed(10, 8),
    to_signed(8, 8),
    to_signed(8, 8),
    to_signed(9, 8),
    to_signed(10, 8),
    to_signed(10, 8),
    to_signed(10, 8),
    to_signed(12, 8),
    to_signed(14, 8),
    to_signed(16, 8),
    to_signed(16, 8),
    to_signed(15, 8),
    to_signed(14, 8),
    to_signed(12, 8),
    to_signed(11, 8),
    to_signed(9, 8),
    to_signed(9, 8),
    to_signed(8, 8),
    to_signed(7, 8),
    to_signed(5, 8),
    to_signed(4, 8),
    to_signed(4, 8),
    to_signed(6, 8),
    to_signed(9, 8),
    to_signed(11, 8),
    to_signed(13, 8),
    to_signed(13, 8),
    to_signed(12, 8),
    to_signed(11, 8),
    to_signed(11, 8),
    to_signed(10, 8),
    to_signed(8, 8),
    to_signed(7, 8),
    to_signed(7, 8),
    to_signed(7, 8),
    to_signed(6, 8),
    to_signed(4, 8),
    to_signed(4, 8),
    to_signed(5, 8),
    to_signed(7, 8),
    to_signed(8, 8),
    to_signed(5, 8),
    to_signed(1, 8),
    to_signed(-1, 8),
    to_signed(1, 8),
    to_signed(4, 8),
    to_signed(6, 8),
    to_signed(6, 8),
    to_signed(8, 8),
    to_signed(12, 8),
    to_signed(13, 8),
    to_signed(10, 8),
    to_signed(6, 8),
    to_signed(3, 8),
    to_signed(2, 8),
    to_signed(2, 8),
    to_signed(3, 8),
    to_signed(3, 8),
    to_signed(3, 8),
    to_signed(2, 8),
    to_signed(3, 8),
    to_signed(3, 8),
    to_signed(1, 8),
    to_signed(-1, 8),
    to_signed(-2, 8),
    to_signed(-2, 8),
    to_signed(0, 8),
    to_signed(2, 8),
    to_signed(5, 8),
    to_signed(4, 8),
    to_signed(1, 8),
    to_signed(-1, 8),
    to_signed(-2, 8),
    to_signed(0, 8),
    to_signed(1, 8),
    to_signed(1, 8),
    to_signed(0, 8),
    to_signed(-1, 8),
    to_signed(-2, 8),
    to_signed(-2, 8),
    to_signed(-3, 8),
    to_signed(-3, 8),
    to_signed(-1, 8),
    to_signed(3, 8),
    to_signed(6, 8),
    to_signed(7, 8),
    to_signed(7, 8),
    to_signed(6, 8),
    to_signed(5, 8),
    to_signed(3, 8),
    to_signed(1, 8),
    to_signed(1, 8),
    to_signed(2, 8),
    to_signed(2, 8),
    to_signed(1, 8),
    to_signed(0, 8),
    to_signed(2, 8),
    to_signed(5, 8),
    to_signed(8, 8),
    to_signed(8, 8),
    to_signed(6, 8),
    to_signed(5, 8),
    to_signed(5, 8),
    to_signed(4, 8),
    to_signed(3, 8),
    to_signed(2, 8),
    to_signed(4, 8),
    to_signed(6, 8),
    to_signed(6, 8),
    to_signed(5, 8),
    to_signed(3, 8),
    to_signed(2, 8),
    to_signed(1, 8),
    to_signed(-2, 8),
    to_signed(-6, 8),
    to_signed(-10, 8),
    to_signed(-10, 8),
    to_signed(-8, 8),
    to_signed(-7, 8),
    to_signed(-6, 8),
    to_signed(-5, 8),
    to_signed(-2, 8),
    to_signed(-1, 8),
    to_signed(-1, 8),
    to_signed(-4, 8),
    to_signed(-6, 8),
    to_signed(-8, 8),
    to_signed(-10, 8),
    to_signed(-12, 8),
    to_signed(-12, 8),
    to_signed(-12, 8),
    to_signed(-12, 8),
    to_signed(-12, 8),
    to_signed(-10, 8),
    to_signed(-7, 8),
    to_signed(-6, 8),
    to_signed(-6, 8),
    to_signed(-8, 8),
    to_signed(-10, 8),
    to_signed(-10, 8),
    to_signed(-9, 8),
    to_signed(-8, 8),
    to_signed(-7, 8),
    to_signed(-7, 8),
    to_signed(-6, 8),
    to_signed(-4, 8),
    to_signed(-3, 8),
    to_signed(-4, 8),
    to_signed(-5, 8),
    to_signed(-4, 8),
    to_signed(-2, 8),
    to_signed(-2, 8),
    to_signed(-5, 8),
    to_signed(-7, 8),
    to_signed(-5, 8),
    to_signed(-3, 8),
    to_signed(-1, 8),
    to_signed(-2, 8),
    to_signed(-3, 8),
    to_signed(-5, 8),
    to_signed(-6, 8),
    to_signed(-7, 8),
    to_signed(-7, 8),
    to_signed(-6, 8),
    to_signed(-6, 8),
    to_signed(-7, 8),
    to_signed(-9, 8),
    to_signed(-11, 8),
    to_signed(-11, 8),
    to_signed(-9, 8),
    to_signed(-6, 8),
    to_signed(-2, 8),
    to_signed(1, 8),
    to_signed(2, 8),
    to_signed(0, 8),
    to_signed(-1, 8),
    to_signed(0, 8),
    to_signed(-1, 8),
    to_signed(-2, 8),
    to_signed(-2, 8),
    to_signed(-1, 8),
    to_signed(-1, 8),
    to_signed(-3, 8),
    to_signed(-6, 8),
    to_signed(-9, 8),
    to_signed(-10, 8),
    to_signed(-11, 8),
    to_signed(-11, 8),
    to_signed(-12, 8),
    to_signed(-14, 8),
    to_signed(-16, 8),
    to_signed(-17, 8),
    to_signed(-15, 8),
    to_signed(-11, 8),
    to_signed(-7, 8),
    to_signed(-3, 8),
    to_signed(-2, 8),
    to_signed(-5, 8),
    to_signed(-10, 8),
    to_signed(-14, 8),
    to_signed(-16, 8),
    to_signed(-16, 8),
    to_signed(-14, 8),
    to_signed(-14, 8),
    to_signed(-15, 8),
    to_signed(-14, 8),
    to_signed(-11, 8),
    to_signed(-9, 8),
    to_signed(-6, 8),
    to_signed(-2, 8),
    to_signed(-1, 8),
    to_signed(-1, 8),
    to_signed(-2, 8),
    to_signed(-4, 8),
    to_signed(-5, 8),
    to_signed(-6, 8),
    to_signed(-4, 8),
    to_signed(-1, 8),
    to_signed(1, 8),
    to_signed(2, 8),
    to_signed(4, 8),
    to_signed(3, 8),
    to_signed(2, 8),
    to_signed(1, 8),
    to_signed(1, 8),
    to_signed(1, 8),
    to_signed(2, 8),
    to_signed(2, 8),
    to_signed(1, 8),
    to_signed(2, 8),
    to_signed(5, 8),
    to_signed(7, 8),
    to_signed(7, 8),
    to_signed(5, 8),
    to_signed(3, 8),
    to_signed(2, 8),
    to_signed(0, 8),
    to_signed(-2, 8),
    to_signed(-2, 8),
    to_signed(0, 8),
    to_signed(1, 8),
    to_signed(-1, 8),
    to_signed(-3, 8),
    to_signed(-5, 8),
    to_signed(-5, 8),
    to_signed(-4, 8),
    to_signed(-3, 8),
    to_signed(-2, 8),
    to_signed(-2, 8),
    to_signed(-3, 8),
    to_signed(-5, 8),
    to_signed(-7, 8),
    to_signed(-8, 8),
    to_signed(-8, 8),
    to_signed(-9, 8),
    to_signed(-10, 8),
    to_signed(-10, 8),
    to_signed(-11, 8),
    to_signed(-13, 8),
    to_signed(-13, 8),
    to_signed(-12, 8),
    to_signed(-10, 8),
    to_signed(-10, 8),
    to_signed(-10, 8),
    to_signed(-9, 8),
    to_signed(-6, 8),
    to_signed(-1, 8),
    to_signed(3, 8),
    to_signed(4, 8),
    to_signed(6, 8),
    to_signed(7, 8),
    to_signed(5, 8),
    to_signed(3, 8),
    to_signed(0, 8),
    to_signed(-1, 8),
    to_signed(0, 8),
    to_signed(1, 8),
    to_signed(3, 8),
    to_signed(5, 8),
    to_signed(6, 8),
    to_signed(6, 8),
    to_signed(5, 8),
    to_signed(2, 8),
    to_signed(-2, 8),
    to_signed(-4, 8),
    to_signed(-2, 8),
    to_signed(3, 8),
    to_signed(5, 8),
    to_signed(4, 8),
    to_signed(2, 8),
    to_signed(3, 8),
    to_signed(6, 8),
    to_signed(8, 8),
    to_signed(7, 8),
    to_signed(4, 8),
    to_signed(2, 8),
    to_signed(0, 8),
    to_signed(0, 8),
    to_signed(2, 8),
    to_signed(6, 8),
    to_signed(8, 8),
    to_signed(8, 8),
    to_signed(4, 8),
    to_signed(3, 8),
    to_signed(4, 8),
    to_signed(6, 8),
    to_signed(5, 8),
    to_signed(4, 8),
    to_signed(5, 8),
    to_signed(6, 8),
    to_signed(5, 8),
    to_signed(3, 8),
    to_signed(3, 8),
    to_signed(5, 8),
    to_signed(7, 8),
    to_signed(6, 8),
    to_signed(3, 8),
    to_signed(0, 8),
    to_signed(0, 8),
    to_signed(2, 8),
    to_signed(5, 8),
    to_signed(8, 8),
    to_signed(8, 8),
    to_signed(6, 8),
    to_signed(5, 8),
    to_signed(6, 8),
    to_signed(8, 8),
    to_signed(9, 8),
    to_signed(9, 8),
    to_signed(7, 8),
    to_signed(4, 8),
    to_signed(2, 8),
    to_signed(-1, 8),
    to_signed(-2, 8),
    to_signed(-2, 8),
    to_signed(-2, 8),
    to_signed(-2, 8),
    to_signed(-1, 8),
    to_signed(2, 8),
    to_signed(6, 8),
    to_signed(8, 8),
    to_signed(7, 8),
    to_signed(5, 8),
    to_signed(4, 8),
    to_signed(3, 8),
    to_signed(-1, 8),
    to_signed(-6, 8),
    to_signed(-7, 8),
    to_signed(-4, 8),
    to_signed(-1, 8),
    to_signed(-1, 8),
    to_signed(0, 8),
    to_signed(3, 8),
    to_signed(6, 8),
    to_signed(6, 8),
    to_signed(2, 8),
    to_signed(-1, 8),
    to_signed(-3, 8),
    to_signed(-4, 8),
    to_signed(-7, 8),
    to_signed(-9, 8),
    to_signed(-10, 8),
    to_signed(-8, 8),
    to_signed(-6, 8),
    to_signed(-3, 8),
    to_signed(-1, 8),
    to_signed(0, 8),
    to_signed(-1, 8),
    to_signed(-4, 8),
    to_signed(-6, 8),
    to_signed(-6, 8),
    to_signed(-5, 8),
    to_signed(-5, 8),
    to_signed(-7, 8),
    to_signed(-11, 8),
    to_signed(-11, 8),
    to_signed(-8, 8),
    to_signed(-7, 8),
    to_signed(-8, 8),
    to_signed(-10, 8),
    to_signed(-10, 8),
    to_signed(-8, 8),
    to_signed(-6, 8),
    to_signed(-6, 8),
    to_signed(-9, 8),
    to_signed(-11, 8),
    to_signed(-11, 8),
    to_signed(-10, 8),
    to_signed(-11, 8),
    to_signed(-12, 8),
    to_signed(-11, 8),
    to_signed(-9, 8),
    to_signed(-7, 8),
    to_signed(-7, 8),
    to_signed(-6, 8),
    to_signed(-5, 8),
    to_signed(-4, 8),
    to_signed(-3, 8),
    to_signed(-3, 8),
    to_signed(-2, 8),
    to_signed(-1, 8),
    to_signed(0, 8),
    to_signed(0, 8),
    to_signed(-3, 8),
    to_signed(-5, 8),
    to_signed(-7, 8),
    to_signed(-8, 8),
    to_signed(-9, 8),
    to_signed(-9, 8),
    to_signed(-6, 8),
    to_signed(-3, 8),
    to_signed(0, 8),
    to_signed(2, 8),
    to_signed(2, 8),
    to_signed(2, 8),
    to_signed(5, 8),
    to_signed(6, 8),
    to_signed(5, 8),
    to_signed(2, 8),
    to_signed(-1, 8),
    to_signed(-2, 8),
    to_signed(-2, 8),
    to_signed(-1, 8),
    to_signed(1, 8),
    to_signed(4, 8),
    to_signed(4, 8),
    to_signed(4, 8),
    to_signed(4, 8),
    to_signed(4, 8),
    to_signed(3, 8),
    to_signed(2, 8),
    to_signed(3, 8),
    to_signed(3, 8),
    to_signed(2, 8),
    to_signed(2, 8),
    to_signed(3, 8),
    to_signed(5, 8),
    to_signed(6, 8),
    to_signed(6, 8),
    to_signed(5, 8),
    to_signed(2, 8),
    to_signed(1, 8),
    to_signed(2, 8),
    to_signed(4, 8),
    to_signed(5, 8),
    to_signed(4, 8),
    to_signed(1, 8),
    to_signed(0, 8),
    to_signed(-1, 8),
    to_signed(-1, 8),
    to_signed(-1, 8),
    to_signed(-2, 8),
    to_signed(-3, 8),
    to_signed(-4, 8),
    to_signed(-4, 8),
    to_signed(-3, 8),
    to_signed(-4, 8),
    to_signed(-4, 8),
    to_signed(-4, 8),
    to_signed(-3, 8),
    to_signed(-3, 8),
    to_signed(-4, 8),
    to_signed(-5, 8),
    to_signed(-4, 8),
    to_signed(-3, 8),
    to_signed(-3, 8),
    to_signed(-3, 8),
    to_signed(-3, 8),
    to_signed(-3, 8),
    to_signed(-2, 8),
    to_signed(-2, 8),
    to_signed(-3, 8),
    to_signed(-3, 8),
    to_signed(-4, 8),
    to_signed(-5, 8),
    to_signed(-6, 8),
    to_signed(-6, 8),
    to_signed(-7, 8),
    to_signed(-9, 8),
    to_signed(-10, 8),
    to_signed(-10, 8),
    to_signed(-9, 8),
    to_signed(-8, 8),
    to_signed(-6, 8),
    to_signed(-3, 8),
    to_signed(0, 8),
    to_signed(1, 8),
    to_signed(1, 8),
    to_signed(0, 8),
    to_signed(0, 8),
    to_signed(-1, 8),
    to_signed(-2, 8),
    to_signed(-3, 8),
    to_signed(-3, 8),
    to_signed(-3, 8),
    to_signed(-3, 8),
    to_signed(-4, 8),
    to_signed(-5, 8),
    to_signed(-3, 8),
    to_signed(0, 8),
    to_signed(1, 8),
    to_signed(2, 8),
    to_signed(2, 8),
    to_signed(2, 8),
    to_signed(3, 8),
    to_signed(4, 8),
    to_signed(6, 8),
    to_signed(5, 8),
    to_signed(3, 8),
    to_signed(4, 8),
    to_signed(6, 8),
    to_signed(8, 8),
    to_signed(8, 8),
    to_signed(6, 8),
    to_signed(5, 8),
    to_signed(5, 8),
    to_signed(4, 8),
    to_signed(2, 8),
    to_signed(2, 8),
    to_signed(3, 8),
    to_signed(5, 8),
    to_signed(8, 8),
    to_signed(8, 8),
    to_signed(7, 8),
    to_signed(7, 8),
    to_signed(7, 8),
    to_signed(6, 8),
    to_signed(6, 8),
    to_signed(7, 8),
    to_signed(8, 8),
    to_signed(8, 8),
    to_signed(7, 8),
    to_signed(8, 8),
    to_signed(10, 8),
    to_signed(11, 8),
    to_signed(11, 8),
    to_signed(9, 8),
    to_signed(7, 8),
    to_signed(7, 8),
    to_signed(10, 8),
    to_signed(14, 8),
    to_signed(15, 8),
    to_signed(14, 8),
    to_signed(12, 8),
    to_signed(12, 8),
    to_signed(14, 8),
    to_signed(17, 8),
    to_signed(20, 8),
    to_signed(20, 8),
    to_signed(18, 8),
    to_signed(16, 8),
    to_signed(14, 8),
    to_signed(12, 8),
    to_signed(12, 8),
    to_signed(13, 8),
    to_signed(14, 8),
    to_signed(12, 8),
    to_signed(11, 8),
    to_signed(11, 8),
    to_signed(13, 8),
    to_signed(14, 8),
    to_signed(13, 8),
    to_signed(12, 8),
    to_signed(11, 8),
    to_signed(8, 8),
    to_signed(6, 8),
    to_signed(5, 8),
    to_signed(4, 8),
    to_signed(4, 8),
    to_signed(4, 8),
    to_signed(2, 8),
    to_signed(-1, 8),
    to_signed(-2, 8),
    to_signed(-3, 8),
    to_signed(-2, 8),
    to_signed(-2, 8),
    to_signed(-1, 8),
    to_signed(1, 8),
    to_signed(3, 8),
    to_signed(4, 8),
    to_signed(4, 8),
    to_signed(2, 8),
    to_signed(-2, 8),
    to_signed(-3, 8),
    to_signed(0, 8),
    to_signed(1, 8),
    to_signed(0, 8),
    to_signed(-2, 8),
    to_signed(-3, 8),
    to_signed(-1, 8),
    to_signed(1, 8),
    to_signed(2, 8),
    to_signed(3, 8),
    to_signed(4, 8),
    to_signed(2, 8),
    to_signed(1, 8),
    to_signed(2, 8),
    to_signed(3, 8),
    to_signed(3, 8),
    to_signed(1, 8),
    to_signed(-1, 8),
    to_signed(-2, 8),
    to_signed(-2, 8),
    to_signed(-2, 8),
    to_signed(-2, 8),
    to_signed(-1, 8),
    to_signed(2, 8),
    to_signed(5, 8),
    to_signed(5, 8),
    to_signed(3, 8),
    to_signed(2, 8),
    to_signed(3, 8),
    to_signed(3, 8),
    to_signed(2, 8),
    to_signed(0, 8),
    to_signed(-1, 8),
    to_signed(0, 8),
    to_signed(0, 8),
    to_signed(3, 8),
    to_signed(7, 8),
    to_signed(8, 8),
    to_signed(7, 8),
    to_signed(5, 8),
    to_signed(4, 8),
    to_signed(3, 8),
    to_signed(3, 8),
    to_signed(3, 8),
    to_signed(3, 8),
    to_signed(1, 8),
    to_signed(0, 8),
    to_signed(0, 8),
    to_signed(1, 8),
    to_signed(1, 8),
    to_signed(-1, 8),
    to_signed(-1, 8),
    to_signed(1, 8),
    to_signed(3, 8),
    to_signed(2, 8),
    to_signed(-2, 8),
    to_signed(-2, 8),
    to_signed(-1, 8),
    to_signed(-2, 8),
    to_signed(-5, 8),
    to_signed(-5, 8),
    to_signed(-2, 8),
    to_signed(0, 8),
    to_signed(-1, 8),
    to_signed(-2, 8),
    to_signed(-3, 8),
    to_signed(-2, 8),
    to_signed(0, 8),
    to_signed(1, 8),
    to_signed(0, 8),
    to_signed(0, 8),
    to_signed(-1, 8),
    to_signed(0, 8),
    to_signed(1, 8),
    to_signed(3, 8),
    to_signed(5, 8),
    to_signed(6, 8),
    to_signed(3, 8),
    to_signed(-1, 8),
    to_signed(0, 8),
    to_signed(2, 8),
    to_signed(3, 8),
    to_signed(2, 8),
    to_signed(2, 8),
    to_signed(2, 8),
    to_signed(2, 8),
    to_signed(3, 8),
    to_signed(3, 8),
    to_signed(0, 8),
    to_signed(-2, 8),
    to_signed(-3, 8),
    to_signed(-2, 8),
    to_signed(-1, 8),
    to_signed(-1, 8),
    to_signed(-1, 8),
    to_signed(0, 8),
    to_signed(3, 8),
    to_signed(3, 8),
    to_signed(2, 8),
    to_signed(1, 8),
    to_signed(2, 8),
    to_signed(3, 8),
    to_signed(5, 8),
    to_signed(7, 8),
    to_signed(7, 8),
    to_signed(6, 8),
    to_signed(3, 8),
    to_signed(0, 8),
    to_signed(-1, 8),
    to_signed(1, 8),
    to_signed(2, 8),
    to_signed(2, 8),
    to_signed(1, 8),
    to_signed(-1, 8),
    to_signed(-1, 8),
    to_signed(-2, 8),
    to_signed(-2, 8),
    to_signed(-2, 8),
    to_signed(-3, 8),
    to_signed(-3, 8),
    to_signed(-2, 8),
    to_signed(-3, 8),
    to_signed(-4, 8),
    to_signed(-8, 8),
    to_signed(-10, 8),
    to_signed(-8, 8),
    to_signed(-5, 8),
    to_signed(-5, 8),
    to_signed(-6, 8),
    to_signed(-7, 8),
    to_signed(-8, 8),
    to_signed(-10, 8),
    to_signed(-12, 8),
    to_signed(-13, 8),
    to_signed(-11, 8),
    to_signed(-8, 8),
    to_signed(-9, 8),
    to_signed(-12, 8),
    to_signed(-15, 8),
    to_signed(-15, 8),
    to_signed(-13, 8),
    to_signed(-10, 8),
    to_signed(-9, 8),
    to_signed(-10, 8),
    to_signed(-11, 8),
    to_signed(-10, 8),
    to_signed(-7, 8),
    to_signed(-3, 8),
    to_signed(0, 8),
    to_signed(-1, 8),
    to_signed(-6, 8),
    to_signed(-9, 8),
    to_signed(-10, 8),
    to_signed(-11, 8),
    to_signed(-12, 8),
    to_signed(-11, 8),
    to_signed(-7, 8),
    to_signed(-6, 8),
    to_signed(-8, 8),
    to_signed(-11, 8),
    to_signed(-11, 8),
    to_signed(-8, 8),
    to_signed(-5, 8),
    to_signed(-5, 8),
    to_signed(-4, 8),
    to_signed(-4, 8),
    to_signed(-6, 8),
    to_signed(-8, 8),
    to_signed(-7, 8),
    to_signed(-5, 8),
    to_signed(-3, 8),
    to_signed(-4, 8),
    to_signed(-6, 8),
    to_signed(-8, 8),
    to_signed(-6, 8),
    to_signed(-3, 8),
    to_signed(-1, 8),
    to_signed(0, 8),
    to_signed(-1, 8),
    to_signed(-3, 8),
    to_signed(-4, 8),
    to_signed(-4, 8),
    to_signed(-5, 8),
    to_signed(-5, 8),
    to_signed(-4, 8),
    to_signed(-4, 8),
    to_signed(-2, 8),
    to_signed(-1, 8),
    to_signed(-1, 8),
    to_signed(-2, 8),
    to_signed(-2, 8),
    to_signed(0, 8),
    to_signed(0, 8),
    to_signed(-2, 8),
    to_signed(-4, 8),
    to_signed(-4, 8),
    to_signed(-3, 8),
    to_signed(-3, 8),
    to_signed(0, 8),
    to_signed(0, 8),
    to_signed(-3, 8),
    to_signed(-7, 8),
    to_signed(-8, 8),
    to_signed(-7, 8),
    to_signed(-5, 8),
    to_signed(-3, 8),
    to_signed(0, 8),
    to_signed(2, 8),
    to_signed(0, 8),
    to_signed(-3, 8),
    to_signed(-5, 8),
    to_signed(-5, 8),
    to_signed(-2, 8),
    to_signed(0, 8),
    to_signed(-1, 8),
    to_signed(-4, 8),
    to_signed(-6, 8),
    to_signed(-5, 8),
    to_signed(-5, 8),
    to_signed(-5, 8),
    to_signed(-6, 8),
    to_signed(-6, 8),
    to_signed(-7, 8),
    to_signed(-9, 8),
    to_signed(-11, 8),
    to_signed(-12, 8),
    to_signed(-10, 8),
    to_signed(-9, 8),
    to_signed(-8, 8),
    to_signed(-8, 8),
    to_signed(-9, 8),
    to_signed(-8, 8),
    to_signed(-5, 8),
    to_signed(-3, 8),
    to_signed(-4, 8),
    to_signed(-4, 8),
    to_signed(-2, 8),
    to_signed(0, 8),
    to_signed(3, 8),
    to_signed(5, 8),
    to_signed(3, 8),
    to_signed(1, 8),
    to_signed(2, 8),
    to_signed(4, 8),
    to_signed(4, 8),
    to_signed(4, 8),
    to_signed(4, 8),
    to_signed(7, 8),
    to_signed(9, 8),
    to_signed(10, 8),
    to_signed(9, 8),
    to_signed(8, 8),
    to_signed(7, 8),
    to_signed(6, 8),
    to_signed(5, 8),
    to_signed(5, 8),
    to_signed(6, 8),
    to_signed(7, 8),
    to_signed(7, 8),
    to_signed(6, 8),
    to_signed(3, 8),
    to_signed(2, 8),
    to_signed(2, 8),
    to_signed(3, 8),
    to_signed(3, 8),
    to_signed(2, 8),
    to_signed(1, 8),
    to_signed(0, 8),
    to_signed(1, 8),
    to_signed(0, 8),
    to_signed(-3, 8),
    to_signed(-3, 8),
    to_signed(-1, 8),
    to_signed(0, 8),
    to_signed(-2, 8),
    to_signed(-5, 8),
    to_signed(-7, 8),
    to_signed(-6, 8),
    to_signed(-6, 8),
    to_signed(-6, 8),
    to_signed(-7, 8),
    to_signed(-7, 8),
    to_signed(-9, 8),
    to_signed(-11, 8),
    to_signed(-11, 8),
    to_signed(-9, 8),
    to_signed(-9, 8),
    to_signed(-9, 8),
    to_signed(-7, 8),
    to_signed(-5, 8),
    to_signed(-4, 8),
    to_signed(-4, 8),
    to_signed(-4, 8),
    to_signed(-5, 8),
    to_signed(-4, 8),
    to_signed(-3, 8),
    to_signed(-4, 8),
    to_signed(-5, 8),
    to_signed(-4, 8),
    to_signed(-2, 8),
    to_signed(-1, 8),
    to_signed(-1, 8),
    to_signed(-2, 8),
    to_signed(-3, 8),
    to_signed(-3, 8),
    to_signed(-4, 8),
    to_signed(-3, 8),
    to_signed(-2, 8),
    to_signed(0, 8),
    to_signed(-1, 8),
    to_signed(-1, 8),
    to_signed(-3, 8),
    to_signed(-6, 8),
    to_signed(-9, 8),
    to_signed(-10, 8),
    to_signed(-10, 8),
    to_signed(-9, 8),
    to_signed(-9, 8),
    to_signed(-8, 8),
    to_signed(-7, 8),
    to_signed(-5, 8),
    to_signed(-4, 8),
    to_signed(-2, 8),
    to_signed(-1, 8),
    to_signed(-1, 8),
    to_signed(-3, 8),
    to_signed(-6, 8),
    to_signed(-7, 8),
    to_signed(-7, 8),
    to_signed(-7, 8),
    to_signed(-7, 8),
    to_signed(-7, 8),
    to_signed(-6, 8),
    to_signed(-5, 8),
    to_signed(-5, 8),
    to_signed(-6, 8),
    to_signed(-6, 8),
    to_signed(-5, 8),
    to_signed(-4, 8),
    to_signed(-1, 8),
    to_signed(3, 8),
    to_signed(4, 8),
    to_signed(1, 8),
    to_signed(1, 8),
    to_signed(5, 8),
    to_signed(8, 8),
    to_signed(6, 8),
    to_signed(2, 8),
    to_signed(1, 8),
    to_signed(3, 8),
    to_signed(6, 8),
    to_signed(7, 8),
    to_signed(7, 8),
    to_signed(6, 8),
    to_signed(4, 8),
    to_signed(2, 8),
    to_signed(-2, 8),
    to_signed(-4, 8),
    to_signed(-2, 8),
    to_signed(2, 8),
    to_signed(5, 8),
    to_signed(5, 8),
    to_signed(5, 8),
    to_signed(6, 8),
    to_signed(9, 8),
    to_signed(11, 8),
    to_signed(13, 8),
    to_signed(12, 8),
    to_signed(10, 8),
    to_signed(7, 8),
    to_signed(5, 8),
    to_signed(4, 8),
    to_signed(5, 8),
    to_signed(6, 8),
    to_signed(6, 8),
    to_signed(5, 8),
    to_signed(5, 8),
    to_signed(5, 8),
    to_signed(4, 8),
    to_signed(2, 8),
    to_signed(2, 8),
    to_signed(4, 8),
    to_signed(5, 8),
    to_signed(6, 8),
    to_signed(6, 8),
    to_signed(5, 8),
    to_signed(3, 8),
    to_signed(1, 8),
    to_signed(0, 8),
    to_signed(0, 8),
    to_signed(0, 8),
    to_signed(0, 8),
    to_signed(1, 8),
    to_signed(1, 8),
    to_signed(-1, 8),
    to_signed(-4, 8),
    to_signed(-7, 8),
    to_signed(-10, 8),
    to_signed(-11, 8),
    to_signed(-11, 8),
    to_signed(-12, 8),
    to_signed(-15, 8),
    to_signed(-17, 8),
    to_signed(-18, 8),
    to_signed(-19, 8),
    to_signed(-18, 8),
    to_signed(-18, 8),
    to_signed(-19, 8),
    to_signed(-19, 8),
    to_signed(-18, 8),
    to_signed(-16, 8),
    to_signed(-16, 8),
    to_signed(-16, 8),
    to_signed(-16, 8),
    to_signed(-13, 8),
    to_signed(-10, 8),
    to_signed(-10, 8),
    to_signed(-11, 8),
    to_signed(-10, 8),
    to_signed(-8, 8),
    to_signed(-5, 8),
    to_signed(-3, 8),
    to_signed(1, 8),
    to_signed(6, 8),
    to_signed(9, 8),
    to_signed(9, 8),
    to_signed(9, 8),
    to_signed(10, 8),
    to_signed(13, 8),
    to_signed(13, 8),
    to_signed(11, 8),
    to_signed(10, 8),
    to_signed(9, 8),
    to_signed(8, 8),
    to_signed(6, 8),
    to_signed(5, 8),
    to_signed(5, 8),
    to_signed(5, 8),
    to_signed(4, 8),
    to_signed(2, 8),
    to_signed(0, 8),
    to_signed(-2, 8),
    to_signed(-2, 8),
    to_signed(-2, 8),
    to_signed(-2, 8),
    to_signed(-3, 8),
    to_signed(-3, 8),
    to_signed(-2, 8),
    to_signed(-1, 8),
    to_signed(0, 8),
    to_signed(3, 8),
    to_signed(7, 8),
    to_signed(8, 8),
    to_signed(6, 8),
    to_signed(5, 8),
    to_signed(7, 8),
    to_signed(9, 8),
    to_signed(8, 8),
    to_signed(7, 8),
    to_signed(6, 8),
    to_signed(6, 8),
    to_signed(7, 8),
    to_signed(7, 8),
    to_signed(8, 8),
    to_signed(8, 8),
    to_signed(8, 8),
    to_signed(7, 8),
    to_signed(8, 8),
    to_signed(9, 8),
    to_signed(9, 8),
    to_signed(9, 8),
    to_signed(8, 8),
    to_signed(7, 8),
    to_signed(7, 8),
    to_signed(8, 8),
    to_signed(9, 8),
    to_signed(9, 8),
    to_signed(9, 8),
    to_signed(8, 8),
    to_signed(7, 8),
    to_signed(6, 8),
    to_signed(5, 8),
    to_signed(5, 8),
    to_signed(5, 8),
    to_signed(5, 8),
    to_signed(4, 8),
    to_signed(5, 8),
    to_signed(6, 8),
    to_signed(6, 8),
    to_signed(7, 8),
    to_signed(9, 8),
    to_signed(10, 8),
    to_signed(9, 8),
    to_signed(9, 8),
    to_signed(9, 8),
    to_signed(8, 8),
    to_signed(6, 8),
    to_signed(4, 8),
    to_signed(4, 8),
    to_signed(4, 8),
    to_signed(3, 8),
    to_signed(0, 8),
    to_signed(-4, 8),
    to_signed(-6, 8),
    to_signed(-6, 8),
    to_signed(-5, 8),
    to_signed(-4, 8),
    to_signed(-4, 8),
    to_signed(-5, 8),
    to_signed(-5, 8),
    to_signed(-4, 8),
    to_signed(-3, 8),
    to_signed(-6, 8),
    to_signed(-8, 8),
    to_signed(-8, 8),
    to_signed(-7, 8),
    to_signed(-8, 8),
    to_signed(-10, 8),
    to_signed(-11, 8),
    to_signed(-10, 8),
    to_signed(-10, 8),
    to_signed(-10, 8),
    to_signed(-10, 8),
    to_signed(-11, 8),
    to_signed(-11, 8),
    to_signed(-9, 8),
    to_signed(-8, 8),
    to_signed(-9, 8),
    to_signed(-10, 8),
    to_signed(-9, 8),
    to_signed(-9, 8),
    to_signed(-11, 8),
    to_signed(-13, 8),
    to_signed(-12, 8),
    to_signed(-11, 8),
    to_signed(-12, 8),
    to_signed(-12, 8),
    to_signed(-10, 8),
    to_signed(-7, 8),
    to_signed(-5, 8),
    to_signed(-5, 8),
    to_signed(-7, 8),
    to_signed(-9, 8),
    to_signed(-10, 8),
    to_signed(-11, 8),
    to_signed(-13, 8),
    to_signed(-16, 8),
    to_signed(-17, 8),
    to_signed(-17, 8),
    to_signed(-18, 8),
    to_signed(-22, 8),
    to_signed(-23, 8),
    to_signed(-21, 8),
    to_signed(-18, 8),
    to_signed(-16, 8),
    to_signed(-15, 8),
    to_signed(-14, 8),
    to_signed(-14, 8),
    to_signed(-15, 8),
    to_signed(-15, 8),
    to_signed(-15, 8),
    to_signed(-16, 8),
    to_signed(-16, 8),
    to_signed(-16, 8),
    to_signed(-16, 8),
    to_signed(-16, 8),
    to_signed(-15, 8),
    to_signed(-15, 8),
    to_signed(-16, 8),
    to_signed(-19, 8),
    to_signed(-22, 8),
    to_signed(-21, 8),
    to_signed(-18, 8),
    to_signed(-17, 8),
    to_signed(-15, 8),
    to_signed(-12, 8),
    to_signed(-10, 8),
    to_signed(-10, 8),
    to_signed(-10, 8),
    to_signed(-9, 8),
    to_signed(-6, 8),
    to_signed(-2, 8),
    to_signed(0, 8),
    to_signed(1, 8),
    to_signed(1, 8),
    to_signed(3, 8),
    to_signed(4, 8),
    to_signed(4, 8),
    to_signed(2, 8),
    to_signed(0, 8),
    to_signed(1, 8),
    to_signed(1, 8),
    to_signed(1, 8),
    to_signed(0, 8),
    to_signed(0, 8),
    to_signed(1, 8),
    to_signed(2, 8),
    to_signed(3, 8),
    to_signed(3, 8),
    to_signed(5, 8),
    to_signed(7, 8),
    to_signed(8, 8),
    to_signed(7, 8),
    to_signed(4, 8),
    to_signed(3, 8),
    to_signed(4, 8),
    to_signed(6, 8),
    to_signed(8, 8),
    to_signed(8, 8),
    to_signed(7, 8),
    to_signed(6, 8),
    to_signed(4, 8),
    to_signed(2, 8),
    to_signed(1, 8),
    to_signed(1, 8),
    to_signed(0, 8),
    to_signed(-2, 8),
    to_signed(-2, 8),
    to_signed(-2, 8),
    to_signed(-2, 8),
    to_signed(-4, 8),
    to_signed(-4, 8),
    to_signed(-4, 8),
    to_signed(-6, 8),
    to_signed(-10, 8),
    to_signed(-14, 8),
    to_signed(-14, 8),
    to_signed(-10, 8),
    to_signed(-6, 8),
    to_signed(-5, 8),
    to_signed(-4, 8),
    to_signed(-2, 8),
    to_signed(1, 8),
    to_signed(2, 8),
    to_signed(1, 8),
    to_signed(-2, 8),
    to_signed(-2, 8),
    to_signed(-1, 8),
    to_signed(-2, 8),
    to_signed(-3, 8),
    to_signed(-3, 8),
    to_signed(-1, 8),
    to_signed(0, 8),
    to_signed(0, 8),
    to_signed(1, 8),
    to_signed(4, 8),
    to_signed(7, 8),
    to_signed(8, 8),
    to_signed(7, 8),
    to_signed(6, 8),
    to_signed(8, 8),
    to_signed(10, 8),
    to_signed(12, 8),
    to_signed(11, 8),
    to_signed(7, 8),
    to_signed(3, 8),
    to_signed(1, 8),
    to_signed(-1, 8),
    to_signed(-2, 8),
    to_signed(-3, 8),
    to_signed(-1, 8),
    to_signed(2, 8),
    to_signed(2, 8),
    to_signed(1, 8),
    to_signed(2, 8),
    to_signed(6, 8),
    to_signed(9, 8),
    to_signed(9, 8),
    to_signed(7, 8),
    to_signed(5, 8),
    to_signed(5, 8),
    to_signed(6, 8),
    to_signed(5, 8),
    to_signed(4, 8),
    to_signed(5, 8),
    to_signed(5, 8),
    to_signed(4, 8),
    to_signed(2, 8),
    to_signed(1, 8),
    to_signed(0, 8),
    to_signed(1, 8),
    to_signed(2, 8),
    to_signed(3, 8),
    to_signed(3, 8),
    to_signed(2, 8),
    to_signed(2, 8),
    to_signed(2, 8),
    to_signed(3, 8),
    to_signed(3, 8),
    to_signed(2, 8),
    to_signed(1, 8),
    to_signed(0, 8),
    to_signed(0, 8),
    to_signed(2, 8),
    to_signed(3, 8),
    to_signed(4, 8),
    to_signed(5, 8),
    to_signed(5, 8),
    to_signed(5, 8),
    to_signed(5, 8),
    to_signed(4, 8),
    to_signed(1, 8),
    to_signed(-1, 8),
    to_signed(0, 8),
    to_signed(5, 8),
    to_signed(8, 8),
    to_signed(9, 8),
    to_signed(11, 8),
    to_signed(14, 8),
    to_signed(16, 8),
    to_signed(15, 8),
    to_signed(13, 8),
    to_signed(13, 8),
    to_signed(13, 8),
    to_signed(14, 8),
    to_signed(15, 8),
    to_signed(15, 8),
    to_signed(15, 8),
    to_signed(14, 8),
    to_signed(14, 8),
    to_signed(13, 8),
    to_signed(10, 8),
    to_signed(8, 8),
    to_signed(8, 8),
    to_signed(9, 8),
    to_signed(10, 8),
    to_signed(11, 8),
    to_signed(10, 8),
    to_signed(8, 8),
    to_signed(8, 8),
    to_signed(9, 8),
    to_signed(11, 8),
    to_signed(11, 8),
    to_signed(12, 8),
    to_signed(13, 8),
    to_signed(13, 8),
    to_signed(10, 8),
    to_signed(8, 8),
    to_signed(7, 8),
    to_signed(7, 8),
    to_signed(6, 8),
    to_signed(4, 8),
    to_signed(3, 8),
    to_signed(2, 8),
    to_signed(1, 8),
    to_signed(1, 8),
    to_signed(2, 8),
    to_signed(3, 8),
    to_signed(3, 8),
    to_signed(2, 8),
    to_signed(1, 8),
    to_signed(1, 8),
    to_signed(0, 8),
    to_signed(-1, 8),
    to_signed(-1, 8),
    to_signed(0, 8),
    to_signed(2, 8),
    to_signed(2, 8),
    to_signed(3, 8),
    to_signed(4, 8),
    to_signed(2, 8),
    to_signed(0, 8),
    to_signed(-1, 8),
    to_signed(0, 8),
    to_signed(0, 8),
    to_signed(-2, 8),
    to_signed(-3, 8),
    to_signed(-4, 8),
    to_signed(-4, 8),
    to_signed(-4, 8),
    to_signed(-2, 8),
    to_signed(-1, 8),
    to_signed(-1, 8),
    to_signed(-1, 8),
    to_signed(1, 8),
    to_signed(2, 8),
    to_signed(3, 8),
    to_signed(5, 8),
    to_signed(6, 8),
    to_signed(6, 8),
    to_signed(3, 8),
    to_signed(0, 8),
    to_signed(-1, 8),
    to_signed(-3, 8),
    to_signed(-4, 8),
    to_signed(-4, 8),
    to_signed(-2, 8),
    to_signed(-2, 8),
    to_signed(-3, 8),
    to_signed(-3, 8),
    to_signed(-3, 8),
    to_signed(-2, 8),
    to_signed(-2, 8),
    to_signed(-3, 8),
    to_signed(-4, 8),
    to_signed(-3, 8),
    to_signed(1, 8),
    to_signed(4, 8),
    to_signed(6, 8),
    to_signed(6, 8),
    to_signed(6, 8),
    to_signed(7, 8),
    to_signed(5, 8),
    to_signed(3, 8),
    to_signed(3, 8),
    to_signed(5, 8),
    to_signed(6, 8),
    to_signed(6, 8),
    to_signed(6, 8),
    to_signed(6, 8),
    to_signed(4, 8),
    to_signed(2, 8),
    to_signed(1, 8),
    to_signed(2, 8),
    to_signed(1, 8),
    to_signed(1, 8),
    to_signed(2, 8),
    to_signed(6, 8),
    to_signed(7, 8),
    to_signed(6, 8),
    to_signed(4, 8),
    to_signed(4, 8),
    to_signed(3, 8),
    to_signed(3, 8),
    to_signed(3, 8),
    to_signed(3, 8),
    to_signed(2, 8),
    to_signed(2, 8),
    to_signed(3, 8),
    to_signed(2, 8),
    to_signed(0, 8),
    to_signed(0, 8),
    to_signed(0, 8),
    to_signed(-2, 8),
    to_signed(-5, 8),
    to_signed(-6, 8),
    to_signed(-4, 8),
    to_signed(-2, 8),
    to_signed(-4, 8),
    to_signed(-5, 8),
    to_signed(-3, 8),
    to_signed(-1, 8),
    to_signed(0, 8),
    to_signed(-2, 8),
    to_signed(-4, 8),
    to_signed(-4, 8),
    to_signed(-3, 8),
    to_signed(-2, 8),
    to_signed(-2, 8),
    to_signed(-2, 8),
    to_signed(-3, 8),
    to_signed(-3, 8),
    to_signed(-4, 8),
    to_signed(-6, 8),
    to_signed(-7, 8),
    to_signed(-5, 8),
    to_signed(-3, 8),
    to_signed(-4, 8),
    to_signed(-7, 8),
    to_signed(-8, 8),
    to_signed(-6, 8),
    to_signed(-4, 8),
    to_signed(-3, 8),
    to_signed(-2, 8),
    to_signed(-2, 8),
    to_signed(-1, 8),
    to_signed(1, 8),
    to_signed(1, 8),
    to_signed(0, 8),
    to_signed(-1, 8),
    to_signed(0, 8),
    to_signed(2, 8),
    to_signed(1, 8),
    to_signed(1, 8),
    to_signed(2, 8),
    to_signed(3, 8),
    to_signed(3, 8),
    to_signed(1, 8),
    to_signed(1, 8),
    to_signed(3, 8),
    to_signed(3, 8),
    to_signed(1, 8),
    to_signed(1, 8),
    to_signed(1, 8),
    to_signed(1, 8),
    to_signed(2, 8),
    to_signed(4, 8),
    to_signed(5, 8),
    to_signed(5, 8),
    to_signed(4, 8),
    to_signed(4, 8),
    to_signed(2, 8),
    to_signed(1, 8),
    to_signed(0, 8),
    to_signed(0, 8),
    to_signed(-1, 8),
    to_signed(-4, 8),
    to_signed(-6, 8),
    to_signed(-6, 8),
    to_signed(-6, 8),
    to_signed(-7, 8),
    to_signed(-8, 8),
    to_signed(-7, 8),
    to_signed(-7, 8),
    to_signed(-8, 8),
    to_signed(-10, 8),
    to_signed(-9, 8),
    to_signed(-8, 8),
    to_signed(-7, 8),
    to_signed(-7, 8),
    to_signed(-7, 8),
    to_signed(-8, 8),
    to_signed(-7, 8),
    to_signed(-6, 8),
    to_signed(-7, 8),
    to_signed(-8, 8),
    to_signed(-7, 8),
    to_signed(-5, 8),
    to_signed(-4, 8),
    to_signed(-6, 8),
    to_signed(-7, 8),
    to_signed(-6, 8),
    to_signed(-5, 8),
    to_signed(-5, 8),
    to_signed(-5, 8),
    to_signed(-5, 8),
    to_signed(-4, 8),
    to_signed(-3, 8),
    to_signed(-2, 8),
    to_signed(0, 8),
    to_signed(2, 8),
    to_signed(3, 8),
    to_signed(4, 8),
    to_signed(5, 8),
    to_signed(4, 8),
    to_signed(4, 8),
    to_signed(6, 8),
    to_signed(7, 8),
    to_signed(7, 8),
    to_signed(6, 8),
    to_signed(7, 8),
    to_signed(7, 8),
    to_signed(6, 8),
    to_signed(5, 8),
    to_signed(5, 8),
    to_signed(7, 8),
    to_signed(7, 8),
    to_signed(7, 8),
    to_signed(8, 8),
    to_signed(11, 8),
    to_signed(14, 8),
    to_signed(16, 8),
    to_signed(18, 8),
    to_signed(18, 8),
    to_signed(18, 8),
    to_signed(16, 8),
    to_signed(15, 8),
    to_signed(14, 8),
    to_signed(14, 8),
    to_signed(14, 8),
    to_signed(16, 8),
    to_signed(16, 8),
    to_signed(14, 8),
    to_signed(10, 8),
    to_signed(6, 8),
    to_signed(5, 8),
    to_signed(4, 8),
    to_signed(4, 8),
    to_signed(4, 8),
    to_signed(2, 8),
    to_signed(0, 8),
    to_signed(-2, 8),
    to_signed(-2, 8),
    to_signed(-3, 8),
    to_signed(-3, 8),
    to_signed(-2, 8),
    to_signed(0, 8),
    to_signed(-1, 8),
    to_signed(-4, 8),
    to_signed(-5, 8),
    to_signed(-6, 8),
    to_signed(-5, 8),
    to_signed(-5, 8),
    to_signed(-5, 8),
    to_signed(-5, 8),
    to_signed(-7, 8),
    to_signed(-8, 8),
    to_signed(-8, 8),
    to_signed(-8, 8),
    to_signed(-9, 8),
    to_signed(-9, 8),
    to_signed(-8, 8),
    to_signed(-6, 8),
    to_signed(-7, 8),
    to_signed(-8, 8),
    to_signed(-8, 8),
    to_signed(-8, 8),
    to_signed(-7, 8),
    to_signed(-6, 8),
    to_signed(-4, 8),
    to_signed(-3, 8),
    to_signed(-3, 8),
    to_signed(-5, 8),
    to_signed(-6, 8),
    to_signed(-8, 8),
    to_signed(-10, 8),
    to_signed(-12, 8),
    to_signed(-13, 8),
    to_signed(-14, 8),
    to_signed(-16, 8),
    to_signed(-17, 8),
    to_signed(-17, 8),
    to_signed(-17, 8),
    to_signed(-16, 8),
    to_signed(-14, 8),
    to_signed(-12, 8),
    to_signed(-11, 8),
    to_signed(-10, 8),
    to_signed(-9, 8),
    to_signed(-9, 8),
    to_signed(-9, 8),
    to_signed(-9, 8),
    to_signed(-8, 8),
    to_signed(-9, 8),
    to_signed(-10, 8),
    to_signed(-11, 8),
    to_signed(-10, 8),
    to_signed(-10, 8),
    to_signed(-12, 8),
    to_signed(-14, 8),
    to_signed(-13, 8),
    to_signed(-12, 8),
    to_signed(-12, 8),
    to_signed(-12, 8),
    to_signed(-13, 8),
    to_signed(-13, 8),
    to_signed(-13, 8),
    to_signed(-14, 8),
    to_signed(-13, 8),
    to_signed(-12, 8),
    to_signed(-10, 8),
    to_signed(-9, 8),
    to_signed(-8, 8),
    to_signed(-7, 8),
    to_signed(-6, 8),
    to_signed(-7, 8),
    to_signed(-8, 8),
    to_signed(-9, 8),
    to_signed(-10, 8),
    to_signed(-11, 8),
    to_signed(-11, 8),
    to_signed(-11, 8),
    to_signed(-11, 8),
    to_signed(-11, 8),
    to_signed(-9, 8),
    to_signed(-7, 8),
    to_signed(-7, 8),
    to_signed(-7, 8),
    to_signed(-8, 8),
    to_signed(-7, 8),
    to_signed(-5, 8),
    to_signed(-3, 8),
    to_signed(-1, 8),
    to_signed(1, 8),
    to_signed(2, 8),
    to_signed(1, 8),
    to_signed(0, 8),
    to_signed(0, 8),
    to_signed(1, 8),
    to_signed(2, 8),
    to_signed(1, 8),
    to_signed(0, 8),
    to_signed(0, 8),
    to_signed(-1, 8),
    to_signed(-2, 8),
    to_signed(-1, 8),
    to_signed(-1, 8),
    to_signed(0, 8),
    to_signed(0, 8),
    to_signed(-1, 8),
    to_signed(-1, 8),
    to_signed(0, 8),
    to_signed(0, 8),
    to_signed(2, 8),
    to_signed(3, 8),
    to_signed(4, 8),
    to_signed(5, 8),
    to_signed(4, 8),
    to_signed(3, 8),
    to_signed(2, 8),
    to_signed(3, 8),
    to_signed(3, 8),
    to_signed(3, 8),
    to_signed(3, 8),
    to_signed(3, 8),
    to_signed(2, 8),
    to_signed(2, 8),
    to_signed(2, 8),
    to_signed(4, 8),
    to_signed(3, 8),
    to_signed(2, 8),
    to_signed(2, 8),
    to_signed(3, 8),
    to_signed(4, 8),
    to_signed(5, 8),
    to_signed(6, 8),
    to_signed(7, 8),
    to_signed(9, 8),
    to_signed(8, 8),
    to_signed(5, 8),
    to_signed(4, 8),
    to_signed(4, 8),
    to_signed(4, 8),
    to_signed(4, 8),
    to_signed(4, 8),
    to_signed(5, 8),
    to_signed(5, 8),
    to_signed(4, 8),
    to_signed(3, 8),
    to_signed(2, 8),
    to_signed(3, 8),
    to_signed(4, 8),
    to_signed(5, 8),
    to_signed(5, 8),
    to_signed(4, 8),
    to_signed(4, 8),
    to_signed(4, 8),
    to_signed(4, 8),
    to_signed(4, 8),
    to_signed(6, 8),
    to_signed(7, 8),
    to_signed(8, 8),
    to_signed(6, 8),
    to_signed(4, 8),
    to_signed(2, 8),
    to_signed(1, 8),
    to_signed(2, 8),
    to_signed(3, 8),
    to_signed(4, 8),
    to_signed(2, 8),
    to_signed(1, 8),
    to_signed(-1, 8),
    to_signed(-2, 8),
    to_signed(-3, 8),
    to_signed(-3, 8),
    to_signed(-2, 8),
    to_signed(-1, 8),
    to_signed(0, 8),
    to_signed(1, 8),
    to_signed(2, 8),
    to_signed(3, 8),
    to_signed(3, 8),
    to_signed(3, 8),
    to_signed(3, 8),
    to_signed(4, 8),
    to_signed(4, 8),
    to_signed(5, 8),
    to_signed(5, 8),
    to_signed(6, 8),
    to_signed(6, 8),
    to_signed(4, 8),
    to_signed(4, 8),
    to_signed(4, 8),
    to_signed(6, 8),
    to_signed(7, 8),
    to_signed(7, 8),
    to_signed(7, 8),
    to_signed(8, 8),
    to_signed(10, 8),
    to_signed(11, 8),
    to_signed(12, 8),
    to_signed(13, 8),
    to_signed(13, 8),
    to_signed(13, 8),
    to_signed(13, 8),
    to_signed(13, 8),
    to_signed(11, 8),
    to_signed(10, 8),
    to_signed(10, 8),
    to_signed(10, 8),
    to_signed(10, 8),
    to_signed(8, 8),
    to_signed(7, 8),
    to_signed(7, 8),
    to_signed(7, 8),
    to_signed(5, 8),
    to_signed(3, 8),
    to_signed(1, 8),
    to_signed(0, 8),
    to_signed(2, 8),
    to_signed(3, 8),
    to_signed(3, 8),
    to_signed(3, 8),
    to_signed(4, 8),
    to_signed(6, 8),
    to_signed(6, 8),
    to_signed(5, 8),
    to_signed(4, 8),
    to_signed(5, 8),
    to_signed(4, 8),
    to_signed(3, 8),
    to_signed(1, 8),
    to_signed(0, 8),
    to_signed(-1, 8),
    to_signed(-2, 8),
    to_signed(-4, 8),
    to_signed(-6, 8),
    to_signed(-8, 8),
    to_signed(-9, 8),
    to_signed(-9, 8),
    to_signed(-7, 8),
    to_signed(-6, 8),
    to_signed(-6, 8),
    to_signed(-7, 8),
    to_signed(-6, 8),
    to_signed(-4, 8),
    to_signed(-1, 8),
    to_signed(-1, 8),
    to_signed(-4, 8),
    to_signed(-6, 8),
    to_signed(-7, 8),
    to_signed(-5, 8),
    to_signed(-4, 8),
    to_signed(-5, 8),
    to_signed(-6, 8),
    to_signed(-5, 8),
    to_signed(-5, 8),
    to_signed(-6, 8),
    to_signed(-8, 8),
    to_signed(-9, 8),
    to_signed(-8, 8),
    to_signed(-7, 8),
    to_signed(-7, 8),
    to_signed(-6, 8),
    to_signed(-5, 8),
    to_signed(-3, 8),
    to_signed(-3, 8),
    to_signed(-4, 8),
    to_signed(-6, 8),
    to_signed(-5, 8),
    to_signed(-2, 8),
    to_signed(1, 8),
    to_signed(1, 8),
    to_signed(-1, 8),
    to_signed(-5, 8),
    to_signed(-6, 8),
    to_signed(-7, 8),
    to_signed(-8, 8),
    to_signed(-10, 8),
    to_signed(-11, 8),
    to_signed(-12, 8),
    to_signed(-11, 8),
    to_signed(-11, 8),
    to_signed(-12, 8),
    to_signed(-12, 8),
    to_signed(-11, 8),
    to_signed(-10, 8),
    to_signed(-10, 8),
    to_signed(-10, 8),
    to_signed(-11, 8),
    to_signed(-12, 8),
    to_signed(-11, 8),
    to_signed(-10, 8),
    to_signed(-9, 8),
    to_signed(-9, 8),
    to_signed(-9, 8),
    to_signed(-10, 8),
    to_signed(-13, 8),
    to_signed(-15, 8),
    to_signed(-16, 8),
    to_signed(-15, 8),
    to_signed(-14, 8),
    to_signed(-13, 8),
    to_signed(-12, 8),
    to_signed(-11, 8),
    to_signed(-12, 8),
    to_signed(-12, 8),
    to_signed(-12, 8),
    to_signed(-11, 8),
    to_signed(-10, 8),
    to_signed(-8, 8),
    to_signed(-6, 8),
    to_signed(-4, 8),
    to_signed(-3, 8),
    to_signed(0, 8),
    to_signed(2, 8),
    to_signed(2, 8),
    to_signed(1, 8),
    to_signed(0, 8),
    to_signed(0, 8),
    to_signed(-1, 8),
    to_signed(-1, 8),
    to_signed(-1, 8),
    to_signed(1, 8),
    to_signed(2, 8),
    to_signed(2, 8),
    to_signed(2, 8),
    to_signed(2, 8),
    to_signed(3, 8),
    to_signed(4, 8),
    to_signed(5, 8),
    to_signed(5, 8),
    to_signed(6, 8),
    to_signed(8, 8),
    to_signed(9, 8),
    to_signed(9, 8),
    to_signed(10, 8),
    to_signed(11, 8),
    to_signed(12, 8),
    to_signed(10, 8),
    to_signed(7, 8),
    to_signed(7, 8),
    to_signed(8, 8),
    to_signed(7, 8),
    to_signed(4, 8),
    to_signed(4, 8),
    to_signed(6, 8),
    to_signed(6, 8),
    to_signed(4, 8),
    to_signed(4, 8),
    to_signed(4, 8),
    to_signed(5, 8),
    to_signed(4, 8),
    to_signed(5, 8),
    to_signed(5, 8),
    to_signed(5, 8),
    to_signed(5, 8),
    to_signed(5, 8),
    to_signed(7, 8),
    to_signed(9, 8),
    to_signed(8, 8),
    to_signed(5, 8),
    to_signed(2, 8),
    to_signed(1, 8),
    to_signed(1, 8),
    to_signed(1, 8),
    to_signed(1, 8),
    to_signed(0, 8),
    to_signed(0, 8),
    to_signed(1, 8),
    to_signed(2, 8),
    to_signed(2, 8),
    to_signed(3, 8),
    to_signed(4, 8),
    to_signed(4, 8),
    to_signed(2, 8),
    to_signed(0, 8),
    to_signed(0, 8),
    to_signed(3, 8),
    to_signed(5, 8),
    to_signed(5, 8),
    to_signed(3, 8),
    to_signed(3, 8),
    to_signed(2, 8),
    to_signed(1, 8),
    to_signed(0, 8),
    to_signed(-3, 8),
    to_signed(-4, 8),
    to_signed(-4, 8),
    to_signed(-5, 8),
    to_signed(-6, 8),
    to_signed(-5, 8),
    to_signed(-2, 8),
    to_signed(-3, 8),
    to_signed(-5, 8),
    to_signed(-5, 8),
    to_signed(-4, 8),
    to_signed(-4, 8),
    to_signed(-6, 8),
    to_signed(-6, 8),
    to_signed(-4, 8),
    to_signed(-2, 8),
    to_signed(0, 8),
    to_signed(1, 8),
    to_signed(0, 8),
    to_signed(-1, 8),
    to_signed(-3, 8),
    to_signed(-4, 8),
    to_signed(-5, 8),
    to_signed(-7, 8),
    to_signed(-7, 8),
    to_signed(-6, 8),
    to_signed(-4, 8),
    to_signed(-5, 8),
    to_signed(-6, 8),
    to_signed(-5, 8),
    to_signed(-4, 8),
    to_signed(-4, 8),
    to_signed(-5, 8),
    to_signed(-7, 8),
    to_signed(-7, 8),
    to_signed(-6, 8),
    to_signed(-4, 8),
    to_signed(-2, 8),
    to_signed(-1, 8),
    to_signed(0, 8),
    to_signed(1, 8),
    to_signed(1, 8),
    to_signed(-1, 8),
    to_signed(-3, 8),
    to_signed(-4, 8),
    to_signed(-3, 8),
    to_signed(-2, 8),
    to_signed(-2, 8),
    to_signed(-2, 8),
    to_signed(-2, 8),
    to_signed(-2, 8),
    to_signed(-2, 8),
    to_signed(-2, 8),
    to_signed(-1, 8),
    to_signed(0, 8),
    to_signed(0, 8),
    to_signed(1, 8),
    to_signed(3, 8),
    to_signed(4, 8),
    to_signed(6, 8),
    to_signed(7, 8),
    to_signed(7, 8),
    to_signed(7, 8),
    to_signed(5, 8),
    to_signed(2, 8),
    to_signed(-1, 8),
    to_signed(-3, 8),
    to_signed(0, 8),
    to_signed(6, 8),
    to_signed(9, 8),
    to_signed(7, 8),
    to_signed(3, 8),
    to_signed(2, 8),
    to_signed(4, 8),
    to_signed(4, 8),
    to_signed(1, 8),
    to_signed(0, 8),
    to_signed(2, 8),
    to_signed(4, 8),
    to_signed(3, 8),
    to_signed(3, 8),
    to_signed(4, 8),
    to_signed(6, 8),
    to_signed(5, 8),
    to_signed(4, 8),
    to_signed(3, 8),
    to_signed(2, 8),
    to_signed(-1, 8),
    to_signed(-3, 8),
    to_signed(-3, 8),
    to_signed(-2, 8),
    to_signed(-2, 8),
    to_signed(-3, 8),
    to_signed(-2, 8),
    to_signed(-2, 8),
    to_signed(-3, 8),
    to_signed(-5, 8),
    to_signed(-5, 8),
    to_signed(-4, 8),
    to_signed(-1, 8),
    to_signed(2, 8),
    to_signed(2, 8),
    to_signed(2, 8),
    to_signed(2, 8),
    to_signed(2, 8),
    to_signed(1, 8),
    to_signed(-1, 8),
    to_signed(-2, 8),
    to_signed(0, 8),
    to_signed(1, 8),
    to_signed(2, 8),
    to_signed(2, 8),
    to_signed(1, 8),
    to_signed(-1, 8),
    to_signed(-4, 8),
    to_signed(-3, 8),
    to_signed(-1, 8),
    to_signed(0, 8),
    to_signed(1, 8),
    to_signed(1, 8),
    to_signed(2, 8),
    to_signed(0, 8),
    to_signed(-1, 8),
    to_signed(1, 8),
    to_signed(5, 8),
    to_signed(7, 8),
    to_signed(6, 8),
    to_signed(5, 8),
    to_signed(6, 8),
    to_signed(6, 8),
    to_signed(6, 8),
    to_signed(4, 8),
    to_signed(3, 8),
    to_signed(2, 8),
    to_signed(2, 8),
    to_signed(1, 8),
    to_signed(1, 8),
    to_signed(2, 8),
    to_signed(2, 8),
    to_signed(3, 8),
    to_signed(4, 8),
    to_signed(4, 8),
    to_signed(5, 8),
    to_signed(5, 8),
    to_signed(5, 8),
    to_signed(5, 8),
    to_signed(6, 8),
    to_signed(7, 8),
    to_signed(9, 8),
    to_signed(9, 8),
    to_signed(7, 8),
    to_signed(4, 8),
    to_signed(1, 8),
    to_signed(-1, 8),
    to_signed(-2, 8),
    to_signed(-1, 8),
    to_signed(1, 8),
    to_signed(2, 8),
    to_signed(3, 8),
    to_signed(1, 8),
    to_signed(0, 8),
    to_signed(0, 8),
    to_signed(2, 8),
    to_signed(4, 8),
    to_signed(6, 8),
    to_signed(6, 8),
    to_signed(8, 8),
    to_signed(10, 8),
    to_signed(13, 8),
    to_signed(13, 8),
    to_signed(14, 8),
    to_signed(15, 8),
    to_signed(16, 8),
    to_signed(16, 8),
    to_signed(13, 8),
    to_signed(10, 8),
    to_signed(10, 8),
    to_signed(12, 8),
    to_signed(13, 8),
    to_signed(13, 8),
    to_signed(13, 8),
    to_signed(12, 8),
    to_signed(13, 8),
    to_signed(13, 8),
    to_signed(13, 8),
    to_signed(13, 8),
    to_signed(13, 8),
    to_signed(14, 8),
    to_signed(16, 8),
    to_signed(16, 8),
    to_signed(15, 8),
    to_signed(15, 8),
    to_signed(15, 8),
    to_signed(14, 8),
    to_signed(13, 8),
    to_signed(12, 8),
    to_signed(11, 8),
    to_signed(11, 8),
    to_signed(10, 8),
    to_signed(9, 8),
    to_signed(9, 8),
    to_signed(9, 8),
    to_signed(9, 8),
    to_signed(7, 8),
    to_signed(7, 8),
    to_signed(7, 8),
    to_signed(7, 8),
    to_signed(6, 8),
    to_signed(4, 8),
    to_signed(4, 8),
    to_signed(4, 8),
    to_signed(5, 8),
    to_signed(6, 8),
    to_signed(8, 8),
    to_signed(9, 8),
    to_signed(7, 8),
    to_signed(5, 8),
    to_signed(3, 8),
    to_signed(2, 8),
    to_signed(2, 8),
    to_signed(0, 8),
    to_signed(-2, 8),
    to_signed(-5, 8),
    to_signed(-7, 8),
    to_signed(-8, 8),
    to_signed(-9, 8),
    to_signed(-9, 8),
    to_signed(-10, 8),
    to_signed(-12, 8),
    to_signed(-13, 8),
    to_signed(-13, 8),
    to_signed(-13, 8),
    to_signed(-12, 8),
    to_signed(-12, 8),
    to_signed(-13, 8),
    to_signed(-12, 8),
    to_signed(-11, 8),
    to_signed(-11, 8),
    to_signed(-13, 8),
    to_signed(-15, 8),
    to_signed(-15, 8),
    to_signed(-13, 8),
    to_signed(-12, 8),
    to_signed(-13, 8),
    to_signed(-14, 8),
    to_signed(-15, 8),
    to_signed(-15, 8),
    to_signed(-15, 8),
    to_signed(-13, 8),
    to_signed(-10, 8),
    to_signed(-10, 8),
    to_signed(-11, 8),
    to_signed(-13, 8),
    to_signed(-12, 8),
    to_signed(-10, 8),
    to_signed(-10, 8),
    to_signed(-10, 8),
    to_signed(-9, 8),
    to_signed(-7, 8),
    to_signed(-5, 8),
    to_signed(-5, 8),
    to_signed(-8, 8),
    to_signed(-10, 8),
    to_signed(-10, 8),
    to_signed(-11, 8),
    to_signed(-13, 8),
    to_signed(-14, 8),
    to_signed(-15, 8),
    to_signed(-14, 8),
    to_signed(-13, 8),
    to_signed(-13, 8),
    to_signed(-13, 8),
    to_signed(-11, 8),
    to_signed(-10, 8),
    to_signed(-9, 8),
    to_signed(-10, 8),
    to_signed(-10, 8),
    to_signed(-9, 8),
    to_signed(-6, 8),
    to_signed(-3, 8),
    to_signed(-2, 8),
    to_signed(-2, 8),
    to_signed(-4, 8),
    to_signed(-5, 8),
    to_signed(-6, 8),
    to_signed(-6, 8),
    to_signed(-7, 8),
    to_signed(-6, 8),
    to_signed(-4, 8),
    to_signed(-2, 8),
    to_signed(-3, 8),
    to_signed(-3, 8),
    to_signed(-4, 8),
    to_signed(-4, 8),
    to_signed(-5, 8),
    to_signed(-5, 8),
    to_signed(-5, 8),
    to_signed(-6, 8),
    to_signed(-6, 8),
    to_signed(-6, 8),
    to_signed(-6, 8),
    to_signed(-4, 8),
    to_signed(-3, 8),
    to_signed(-3, 8),
    to_signed(-3, 8),
    to_signed(-4, 8),
    to_signed(-5, 8),
    to_signed(-7, 8),
    to_signed(-8, 8),
    to_signed(-7, 8),
    to_signed(-6, 8),
    to_signed(-5, 8),
    to_signed(-5, 8),
    to_signed(-6, 8),
    to_signed(-6, 8),
    to_signed(-6, 8),
    to_signed(-7, 8),
    to_signed(-7, 8),
    to_signed(-7, 8),
    to_signed(-6, 8),
    to_signed(-5, 8),
    to_signed(-4, 8),
    to_signed(-3, 8),
    to_signed(0, 8),
    to_signed(3, 8),
    to_signed(2, 8),
    to_signed(-1, 8),
    to_signed(-3, 8),
    to_signed(-4, 8),
    to_signed(-6, 8),
    to_signed(-7, 8),
    to_signed(-6, 8),
    to_signed(-4, 8),
    to_signed(-4, 8),
    to_signed(-5, 8),
    to_signed(-5, 8),
    to_signed(-4, 8),
    to_signed(-3, 8),
    to_signed(-4, 8),
    to_signed(-6, 8),
    to_signed(-6, 8),
    to_signed(-5, 8),
    to_signed(-2, 8),
    to_signed(0, 8),
    to_signed(2, 8),
    to_signed(2, 8),
    to_signed(1, 8),
    to_signed(0, 8),
    to_signed(-3, 8),
    to_signed(-4, 8),
    to_signed(-4, 8),
    to_signed(-3, 8),
    to_signed(-3, 8),
    to_signed(-3, 8),
    to_signed(-3, 8),
    to_signed(-2, 8),
    to_signed(-2, 8),
    to_signed(-3, 8),
    to_signed(-3, 8),
    to_signed(-2, 8),
    to_signed(-3, 8),
    to_signed(-5, 8),
    to_signed(-5, 8),
    to_signed(-3, 8),
    to_signed(-1, 8),
    to_signed(0, 8),
    to_signed(2, 8),
    to_signed(4, 8),
    to_signed(4, 8),
    to_signed(1, 8),
    to_signed(-2, 8),
    to_signed(-3, 8),
    to_signed(-2, 8),
    to_signed(-2, 8),
    to_signed(-2, 8),
    to_signed(-2, 8),
    to_signed(-2, 8),
    to_signed(-2, 8),
    to_signed(-3, 8),
    to_signed(-4, 8),
    to_signed(-4, 8),
    to_signed(-5, 8),
    to_signed(-4, 8),
    to_signed(-4, 8),
    to_signed(-4, 8),
    to_signed(-3, 8),
    to_signed(-1, 8),
    to_signed(0, 8),
    to_signed(0, 8),
    to_signed(0, 8),
    to_signed(-1, 8),
    to_signed(-4, 8),
    to_signed(-6, 8),
    to_signed(-7, 8),
    to_signed(-6, 8),
    to_signed(-5, 8),
    to_signed(-4, 8),
    to_signed(-3, 8),
    to_signed(-2, 8),
    to_signed(-3, 8),
    to_signed(-4, 8),
    to_signed(-5, 8),
    to_signed(-6, 8),
    to_signed(-7, 8),
    to_signed(-7, 8),
    to_signed(-5, 8),
    to_signed(-5, 8),
    to_signed(-4, 8),
    to_signed(-4, 8),
    to_signed(-3, 8),
    to_signed(-3, 8),
    to_signed(-4, 8),
    to_signed(-5, 8),
    to_signed(-6, 8),
    to_signed(-7, 8),
    to_signed(-7, 8),
    to_signed(-7, 8),
    to_signed(-7, 8),
    to_signed(-7, 8),
    to_signed(-6, 8),
    to_signed(-7, 8),
    to_signed(-9, 8),
    to_signed(-9, 8),
    to_signed(-9, 8),
    to_signed(-9, 8),
    to_signed(-9, 8),
    to_signed(-9, 8),
    to_signed(-7, 8),
    to_signed(-6, 8),
    to_signed(-7, 8),
    to_signed(-6, 8),
    to_signed(-5, 8),
    to_signed(-4, 8),
    to_signed(-4, 8),
    to_signed(-6, 8),
    to_signed(-6, 8),
    to_signed(-5, 8),
    to_signed(-4, 8),
    to_signed(-4, 8),
    to_signed(-5, 8),
    to_signed(-5, 8),
    to_signed(-3, 8),
    to_signed(-3, 8),
    to_signed(-5, 8),
    to_signed(-7, 8),
    to_signed(-7, 8),
    to_signed(-6, 8),
    to_signed(-7, 8),
    to_signed(-8, 8),
    to_signed(-7, 8),
    to_signed(-5, 8),
    to_signed(-3, 8),
    to_signed(-3, 8),
    to_signed(-4, 8),
    to_signed(-4, 8),
    to_signed(-5, 8),
    to_signed(-8, 8),
    to_signed(-9, 8),
    to_signed(-9, 8),
    to_signed(-7, 8),
    to_signed(-8, 8),
    to_signed(-9, 8),
    to_signed(-10, 8),
    to_signed(-10, 8),
    to_signed(-10, 8),
    to_signed(-11, 8),
    to_signed(-10, 8),
    to_signed(-9, 8),
    to_signed(-8, 8),
    to_signed(-8, 8),
    to_signed(-9, 8),
    to_signed(-8, 8),
    to_signed(-7, 8),
    to_signed(-6, 8),
    to_signed(-6, 8),
    to_signed(-4, 8),
    to_signed(-2, 8),
    to_signed(0, 8),
    to_signed(1, 8),
    to_signed(2, 8),
    to_signed(3, 8),
    to_signed(3, 8),
    to_signed(3, 8),
    to_signed(4, 8),
    to_signed(5, 8),
    to_signed(5, 8),
    to_signed(5, 8),
    to_signed(7, 8),
    to_signed(9, 8),
    to_signed(10, 8),
    to_signed(9, 8),
    to_signed(10, 8),
    to_signed(11, 8),
    to_signed(11, 8),
    to_signed(12, 8),
    to_signed(12, 8),
    to_signed(12, 8),
    to_signed(12, 8),
    to_signed(12, 8),
    to_signed(13, 8),
    to_signed(13, 8),
    to_signed(13, 8),
    to_signed(11, 8),
    to_signed(9, 8),
    to_signed(8, 8),
    to_signed(8, 8),
    to_signed(10, 8),
    to_signed(10, 8),
    to_signed(9, 8),
    to_signed(8, 8),
    to_signed(9, 8),
    to_signed(8, 8),
    to_signed(8, 8),
    to_signed(7, 8),
    to_signed(7, 8),
    to_signed(6, 8),
    to_signed(5, 8),
    to_signed(4, 8),
    to_signed(5, 8),
    to_signed(6, 8),
    to_signed(6, 8),
    to_signed(6, 8),
    to_signed(5, 8),
    to_signed(4, 8),
    to_signed(2, 8),
    to_signed(0, 8),
    to_signed(-1, 8),
    to_signed(0, 8),
    to_signed(1, 8),
    to_signed(1, 8),
    to_signed(1, 8),
    to_signed(2, 8),
    to_signed(2, 8),
    to_signed(1, 8),
    to_signed(-1, 8),
    to_signed(0, 8),
    to_signed(1, 8),
    to_signed(1, 8),
    to_signed(2, 8),
    to_signed(3, 8),
    to_signed(4, 8),
    to_signed(5, 8),
    to_signed(5, 8),
    to_signed(6, 8),
    to_signed(5, 8),
    to_signed(3, 8),
    to_signed(3, 8),
    to_signed(3, 8),
    to_signed(3, 8),
    to_signed(3, 8),
    to_signed(4, 8),
    to_signed(5, 8),
    to_signed(5, 8),
    to_signed(5, 8),
    to_signed(4, 8),
    to_signed(3, 8),
    to_signed(2, 8),
    to_signed(3, 8),
    to_signed(3, 8),
    to_signed(3, 8),
    to_signed(3, 8),
    to_signed(5, 8),
    to_signed(6, 8),
    to_signed(4, 8),
    to_signed(4, 8),
    to_signed(3, 8),
    to_signed(1, 8),
    to_signed(0, 8),
    to_signed(0, 8),
    to_signed(3, 8),
    to_signed(4, 8),
    to_signed(4, 8),
    to_signed(3, 8),
    to_signed(0, 8),
    to_signed(-1, 8),
    to_signed(-1, 8),
    to_signed(0, 8),
    to_signed(-2, 8),
    to_signed(-3, 8),
    to_signed(-2, 8),
    to_signed(0, 8),
    to_signed(1, 8),
    to_signed(1, 8),
    to_signed(0, 8),
    to_signed(-1, 8),
    to_signed(0, 8),
    to_signed(1, 8),
    to_signed(2, 8),
    to_signed(1, 8),
    to_signed(0, 8),
    to_signed(0, 8),
    to_signed(0, 8),
    to_signed(0, 8),
    to_signed(0, 8),
    to_signed(0, 8),
    to_signed(1, 8),
    to_signed(3, 8),
    to_signed(4, 8),
    to_signed(4, 8),
    to_signed(2, 8),
    to_signed(3, 8),
    to_signed(5, 8),
    to_signed(5, 8),
    to_signed(5, 8),
    to_signed(6, 8),
    to_signed(8, 8),
    to_signed(7, 8),
    to_signed(7, 8),
    to_signed(7, 8),
    to_signed(8, 8),
    to_signed(7, 8),
    to_signed(6, 8),
    to_signed(6, 8),
    to_signed(6, 8),
    to_signed(5, 8),
    to_signed(4, 8),
    to_signed(5, 8),
    to_signed(5, 8),
    to_signed(5, 8),
    to_signed(5, 8),
    to_signed(4, 8),
    to_signed(3, 8),
    to_signed(1, 8),
    to_signed(-1, 8),
    to_signed(-1, 8),
    to_signed(0, 8),
    to_signed(0, 8),
    to_signed(0, 8),
    to_signed(0, 8),
    to_signed(0, 8),
    to_signed(0, 8),
    to_signed(-1, 8),
    to_signed(-2, 8),
    to_signed(-2, 8),
    to_signed(-3, 8),
    to_signed(-3, 8),
    to_signed(-1, 8),
    to_signed(1, 8),
    to_signed(2, 8),
    to_signed(1, 8),
    to_signed(1, 8),
    to_signed(1, 8),
    to_signed(1, 8),
    to_signed(1, 8),
    to_signed(2, 8),
    to_signed(3, 8),
    to_signed(2, 8),
    to_signed(2, 8),
    to_signed(3, 8),
    to_signed(3, 8),
    to_signed(3, 8),
    to_signed(3, 8),
    to_signed(4, 8),
    to_signed(5, 8),
    to_signed(5, 8),
    to_signed(5, 8),
    to_signed(5, 8),
    to_signed(6, 8),
    to_signed(6, 8),
    to_signed(6, 8),
    to_signed(5, 8),
    to_signed(5, 8),
    to_signed(6, 8),
    to_signed(6, 8),
    to_signed(7, 8),
    to_signed(8, 8),
    to_signed(8, 8),
    to_signed(7, 8),
    to_signed(7, 8),
    to_signed(8, 8),
    to_signed(8, 8),
    to_signed(7, 8),
    to_signed(6, 8),
    to_signed(5, 8),
    to_signed(6, 8),
    to_signed(7, 8),
    to_signed(7, 8),
    to_signed(7, 8),
    to_signed(6, 8),
    to_signed(5, 8),
    to_signed(4, 8),
    to_signed(2, 8),
    to_signed(1, 8),
    to_signed(1, 8),
    to_signed(2, 8),
    to_signed(3, 8),
    to_signed(4, 8),
    to_signed(3, 8),
    to_signed(2, 8),
    to_signed(0, 8),
    to_signed(0, 8),
    to_signed(0, 8),
    to_signed(0, 8),
    to_signed(0, 8),
    to_signed(0, 8),
    to_signed(-2, 8),
    to_signed(-4, 8),
    to_signed(-4, 8),
    to_signed(-3, 8),
    to_signed(-3, 8),
    to_signed(-5, 8),
    to_signed(-6, 8),
    to_signed(-6, 8),
    to_signed(-4, 8),
    to_signed(-4, 8),
    to_signed(-5, 8),
    to_signed(-6, 8),
    to_signed(-5, 8),
    to_signed(-3, 8),
    to_signed(-1, 8),
    to_signed(-1, 8),
    to_signed(-1, 8),
    to_signed(-2, 8),
    to_signed(-2, 8),
    to_signed(-2, 8),
    to_signed(-1, 8),
    to_signed(0, 8),
    to_signed(2, 8),
    to_signed(2, 8),
    to_signed(3, 8),
    to_signed(3, 8),
    to_signed(3, 8),
    to_signed(3, 8),
    to_signed(2, 8),
    to_signed(2, 8),
    to_signed(2, 8),
    to_signed(3, 8),
    to_signed(3, 8),
    to_signed(3, 8),
    to_signed(3, 8),
    to_signed(4, 8),
    to_signed(4, 8),
    to_signed(4, 8),
    to_signed(3, 8),
    to_signed(2, 8),
    to_signed(1, 8),
    to_signed(-1, 8),
    to_signed(-2, 8),
    to_signed(-2, 8),
    to_signed(-1, 8),
    to_signed(0, 8),
    to_signed(1, 8),
    to_signed(0, 8),
    to_signed(-3, 8),
    to_signed(-4, 8),
    to_signed(-5, 8),
    to_signed(-6, 8),
    to_signed(-6, 8),
    to_signed(-6, 8),
    to_signed(-5, 8),
    to_signed(-4, 8),
    to_signed(-4, 8),
    to_signed(-4, 8),
    to_signed(-5, 8),
    to_signed(-5, 8),
    to_signed(-5, 8),
    to_signed(-5, 8),
    to_signed(-5, 8),
    to_signed(-6, 8),
    to_signed(-5, 8),
    to_signed(-4, 8),
    to_signed(-2, 8),
    to_signed(-2, 8),
    to_signed(-2, 8),
    to_signed(-4, 8),
    to_signed(-6, 8),
    to_signed(-5, 8),
    to_signed(-4, 8),
    to_signed(-4, 8),
    to_signed(-4, 8),
    to_signed(-2, 8),
    to_signed(-1, 8),
    to_signed(-1, 8),
    to_signed(-1, 8),
    to_signed(-1, 8),
    to_signed(0, 8),
    to_signed(0, 8),
    to_signed(0, 8),
    to_signed(0, 8),
    to_signed(0, 8),
    to_signed(-1, 8),
    to_signed(-1, 8),
    to_signed(-1, 8),
    to_signed(0, 8),
    to_signed(-1, 8),
    to_signed(-2, 8),
    to_signed(-2, 8),
    to_signed(-2, 8),
    to_signed(-1, 8),
    to_signed(-2, 8),
    to_signed(-2, 8),
    to_signed(-2, 8),
    to_signed(-1, 8),
    to_signed(1, 8),
    to_signed(1, 8),
    to_signed(2, 8),
    to_signed(4, 8),
    to_signed(5, 8),
    to_signed(6, 8),
    to_signed(6, 8),
    to_signed(6, 8),
    to_signed(6, 8),
    to_signed(5, 8),
    to_signed(3, 8),
    to_signed(3, 8),
    to_signed(4, 8),
    to_signed(6, 8),
    to_signed(6, 8),
    to_signed(5, 8),
    to_signed(2, 8),
    to_signed(2, 8),
    to_signed(2, 8),
    to_signed(2, 8),
    to_signed(1, 8),
    to_signed(0, 8),
    to_signed(-2, 8),
    to_signed(-3, 8),
    to_signed(-4, 8),
    to_signed(-3, 8),
    to_signed(-1, 8),
    to_signed(-1, 8),
    to_signed(-1, 8),
    to_signed(0, 8),
    to_signed(-1, 8),
    to_signed(-4, 8),
    to_signed(-6, 8),
    to_signed(-7, 8),
    to_signed(-6, 8),
    to_signed(-5, 8),
    to_signed(-4, 8),
    to_signed(-3, 8),
    to_signed(-3, 8),
    to_signed(-4, 8),
    to_signed(-4, 8),
    to_signed(-5, 8),
    to_signed(-5, 8),
    to_signed(-6, 8),
    to_signed(-6, 8),
    to_signed(-4, 8),
    to_signed(-3, 8),
    to_signed(-1, 8),
    to_signed(-1, 8),
    to_signed(0, 8),
    to_signed(0, 8),
    to_signed(-1, 8),
    to_signed(-2, 8),
    to_signed(-1, 8),
    to_signed(0, 8),
    to_signed(1, 8),
    to_signed(2, 8),
    to_signed(3, 8),
    to_signed(4, 8),
    to_signed(4, 8),
    to_signed(3, 8),
    to_signed(2, 8),
    to_signed(1, 8),
    to_signed(1, 8),
    to_signed(1, 8),
    to_signed(1, 8),
    to_signed(2, 8),
    to_signed(3, 8),
    to_signed(4, 8),
    to_signed(6, 8),
    to_signed(7, 8),
    to_signed(6, 8),
    to_signed(5, 8),
    to_signed(4, 8),
    to_signed(4, 8),
    to_signed(4, 8),
    to_signed(4, 8),
    to_signed(4, 8),
    to_signed(5, 8),
    to_signed(5, 8),
    to_signed(4, 8),
    to_signed(2, 8),
    to_signed(1, 8),
    to_signed(1, 8),
    to_signed(0, 8),
    to_signed(-1, 8),
    to_signed(0, 8),
    to_signed(2, 8),
    to_signed(3, 8),
    to_signed(3, 8),
    to_signed(1, 8),
    to_signed(0, 8),
    to_signed(0, 8),
    to_signed(1, 8),
    to_signed(1, 8),
    to_signed(3, 8),
    to_signed(5, 8),
    to_signed(5, 8),
    to_signed(3, 8),
    to_signed(0, 8),
    to_signed(-2, 8),
    to_signed(-2, 8),
    to_signed(-2, 8),
    to_signed(-1, 8),
    to_signed(-1, 8),
    to_signed(-1, 8),
    to_signed(0, 8),
    to_signed(-1, 8),
    to_signed(-2, 8),
    to_signed(-3, 8),
    to_signed(-2, 8),
    to_signed(0, 8),
    to_signed(1, 8),
    to_signed(1, 8),
    to_signed(2, 8),
    to_signed(4, 8),
    to_signed(4, 8),
    to_signed(3, 8),
    to_signed(2, 8),
    to_signed(1, 8),
    to_signed(0, 8),
    to_signed(-1, 8),
    to_signed(-1, 8),
    to_signed(0, 8),
    to_signed(0, 8),
    to_signed(-1, 8),
    to_signed(-3, 8),
    to_signed(-5, 8),
    to_signed(-5, 8),
    to_signed(-4, 8),
    to_signed(-4, 8),
    to_signed(-3, 8),
    to_signed(-2, 8),
    to_signed(-1, 8),
    to_signed(-2, 8),
    to_signed(-2, 8),
    to_signed(-2, 8),
    to_signed(-3, 8),
    to_signed(-4, 8),
    to_signed(-5, 8),
    to_signed(-6, 8),
    to_signed(-6, 8),
    to_signed(-5, 8),
    to_signed(-4, 8),
    to_signed(-6, 8),
    to_signed(-9, 8),
    to_signed(-10, 8),
    to_signed(-10, 8),
    to_signed(-9, 8),
    to_signed(-9, 8),
    to_signed(-9, 8),
    to_signed(-7, 8),
    to_signed(-6, 8),
    to_signed(-7, 8),
    to_signed(-9, 8),
    to_signed(-9, 8),
    to_signed(-8, 8),
    to_signed(-8, 8),
    to_signed(-9, 8),
    to_signed(-9, 8),
    to_signed(-9, 8),
    to_signed(-10, 8),
    to_signed(-10, 8),
    to_signed(-10, 8),
    to_signed(-9, 8),
    to_signed(-8, 8),
    to_signed(-9, 8),
    to_signed(-9, 8),
    to_signed(-9, 8),
    to_signed(-10, 8),
    to_signed(-11, 8),
    to_signed(-10, 8),
    to_signed(-10, 8),
    to_signed(-10, 8),
    to_signed(-9, 8),
    to_signed(-9, 8),
    to_signed(-8, 8),
    to_signed(-6, 8),
    to_signed(-5, 8),
    to_signed(-5, 8),
    to_signed(-6, 8),
    to_signed(-7, 8),
    to_signed(-7, 8),
    to_signed(-5, 8),
    to_signed(-5, 8),
    to_signed(-6, 8),
    to_signed(-6, 8),
    to_signed(-6, 8),
    to_signed(-5, 8),
    to_signed(-5, 8),
    to_signed(-6, 8),
    to_signed(-7, 8),
    to_signed(-6, 8),
    to_signed(-6, 8),
    to_signed(-6, 8),
    to_signed(-7, 8),
    to_signed(-7, 8),
    to_signed(-5, 8),
    to_signed(-3, 8),
    to_signed(-2, 8),
    to_signed(-3, 8),
    to_signed(-4, 8),
    to_signed(-6, 8),
    to_signed(-6, 8),
    to_signed(-6, 8),
    to_signed(-5, 8),
    to_signed(-4, 8),
    to_signed(-3, 8),
    to_signed(-2, 8),
    to_signed(-1, 8),
    to_signed(-2, 8),
    to_signed(-3, 8),
    to_signed(-4, 8),
    to_signed(-5, 8),
    to_signed(-6, 8),
    to_signed(-6, 8),
    to_signed(-5, 8),
    to_signed(-4, 8),
    to_signed(-4, 8),
    to_signed(-4, 8),
    to_signed(-3, 8),
    to_signed(-2, 8),
    to_signed(0, 8),
    to_signed(1, 8),
    to_signed(2, 8),
    to_signed(3, 8),
    to_signed(3, 8),
    to_signed(2, 8),
    to_signed(2, 8),
    to_signed(2, 8),
    to_signed(3, 8),
    to_signed(3, 8),
    to_signed(5, 8),
    to_signed(6, 8),
    to_signed(7, 8),
    to_signed(6, 8),
    to_signed(5, 8),
    to_signed(4, 8),
    to_signed(5, 8),
    to_signed(7, 8),
    to_signed(8, 8),
    to_signed(8, 8),
    to_signed(7, 8),
    to_signed(8, 8),
    to_signed(9, 8),
    to_signed(9, 8),
    to_signed(8, 8),
    to_signed(6, 8),
    to_signed(4, 8),
    to_signed(4, 8),
    to_signed(5, 8),
    to_signed(6, 8),
    to_signed(7, 8),
    to_signed(7, 8),
    to_signed(5, 8),
    to_signed(3, 8),
    to_signed(2, 8),
    to_signed(4, 8),
    to_signed(4, 8),
    to_signed(3, 8),
    to_signed(1, 8),
    to_signed(1, 8),
    to_signed(2, 8),
    to_signed(1, 8),
    to_signed(1, 8),
    to_signed(0, 8),
    to_signed(-1, 8),
    to_signed(-2, 8),
    to_signed(-3, 8),
    to_signed(-4, 8),
    to_signed(-5, 8),
    to_signed(-5, 8),
    to_signed(-6, 8),
    to_signed(-6, 8),
    to_signed(-7, 8),
    to_signed(-6, 8),
    to_signed(-6, 8),
    to_signed(-5, 8),
    to_signed(-6, 8),
    to_signed(-8, 8),
    to_signed(-9, 8),
    to_signed(-9, 8),
    to_signed(-10, 8),
    to_signed(-12, 8),
    to_signed(-12, 8),
    to_signed(-11, 8),
    to_signed(-9, 8),
    to_signed(-7, 8),
    to_signed(-7, 8),
    to_signed(-7, 8),
    to_signed(-7, 8),
    to_signed(-7, 8),
    to_signed(-6, 8),
    to_signed(-6, 8),
    to_signed(-6, 8),
    to_signed(-5, 8),
    to_signed(-3, 8),
    to_signed(-1, 8),
    to_signed(0, 8),
    to_signed(-1, 8),
    to_signed(-2, 8),
    to_signed(-2, 8),
    to_signed(-3, 8),
    to_signed(-3, 8),
    to_signed(-4, 8),
    to_signed(-3, 8),
    to_signed(-1, 8),
    to_signed(2, 8),
    to_signed(3, 8),
    to_signed(2, 8),
    to_signed(1, 8),
    to_signed(2, 8),
    to_signed(3, 8),
    to_signed(3, 8),
    to_signed(3, 8),
    to_signed(2, 8),
    to_signed(2, 8),
    to_signed(3, 8),
    to_signed(4, 8),
    to_signed(3, 8),
    to_signed(2, 8),
    to_signed(0, 8),
    to_signed(-1, 8),
    to_signed(-3, 8),
    to_signed(-4, 8),
    to_signed(-4, 8),
    to_signed(-4, 8),
    to_signed(-5, 8),
    to_signed(-4, 8),
    to_signed(-2, 8),
    to_signed(-2, 8),
    to_signed(-2, 8),
    to_signed(-3, 8),
    to_signed(-2, 8),
    to_signed(-3, 8),
    to_signed(-4, 8),
    to_signed(-5, 8),
    to_signed(-5, 8),
    to_signed(-5, 8),
    to_signed(-4, 8),
    to_signed(-4, 8),
    to_signed(-5, 8),
    to_signed(-5, 8),
    to_signed(-7, 8),
    to_signed(-8, 8),
    to_signed(-9, 8),
    to_signed(-9, 8),
    to_signed(-7, 8),
    to_signed(-5, 8),
    to_signed(-6, 8),
    to_signed(-5, 8),
    to_signed(-4, 8),
    to_signed(-3, 8),
    to_signed(-3, 8),
    to_signed(-2, 8),
    to_signed(-1, 8),
    to_signed(-1, 8),
    to_signed(-1, 8),
    to_signed(0, 8),
    to_signed(0, 8),
    to_signed(-1, 8),
    to_signed(-1, 8),
    to_signed(0, 8),
    to_signed(2, 8),
    to_signed(3, 8),
    to_signed(2, 8),
    to_signed(2, 8),
    to_signed(1, 8),
    to_signed(1, 8),
    to_signed(0, 8),
    to_signed(1, 8),
    to_signed(2, 8),
    to_signed(3, 8),
    to_signed(4, 8),
    to_signed(5, 8),
    to_signed(5, 8),
    to_signed(5, 8),
    to_signed(5, 8),
    to_signed(4, 8),
    to_signed(3, 8),
    to_signed(3, 8),
    to_signed(3, 8),
    to_signed(3, 8),
    to_signed(1, 8),
    to_signed(-1, 8),
    to_signed(-2, 8),
    to_signed(-3, 8),
    to_signed(-3, 8),
    to_signed(-4, 8),
    to_signed(-5, 8),
    to_signed(-6, 8),
    to_signed(-6, 8),
    to_signed(-5, 8),
    to_signed(-5, 8),
    to_signed(-5, 8),
    to_signed(-5, 8),
    to_signed(-4, 8),
    to_signed(-4, 8),
    to_signed(-4, 8),
    to_signed(-4, 8),
    to_signed(-5, 8),
    to_signed(-5, 8),
    to_signed(-4, 8),
    to_signed(-5, 8),
    to_signed(-5, 8),
    to_signed(-5, 8),
    to_signed(-2, 8),
    to_signed(-1, 8),
    to_signed(0, 8),
    to_signed(-1, 8),
    to_signed(-1, 8),
    to_signed(-2, 8),
    to_signed(-2, 8),
    to_signed(-1, 8),
    to_signed(0, 8),
    to_signed(1, 8),
    to_signed(3, 8),
    to_signed(4, 8),
    to_signed(5, 8),
    to_signed(6, 8),
    to_signed(7, 8),
    to_signed(6, 8),
    to_signed(6, 8),
    to_signed(7, 8),
    to_signed(8, 8),
    to_signed(9, 8),
    to_signed(9, 8),
    to_signed(10, 8),
    to_signed(11, 8),
    to_signed(11, 8),
    to_signed(10, 8),
    to_signed(9, 8),
    to_signed(7, 8),
    to_signed(5, 8),
    to_signed(4, 8),
    to_signed(5, 8),
    to_signed(6, 8),
    to_signed(8, 8),
    to_signed(8, 8),
    to_signed(7, 8),
    to_signed(7, 8),
    to_signed(7, 8),
    to_signed(6, 8),
    to_signed(5, 8),
    to_signed(4, 8),
    to_signed(4, 8),
    to_signed(4, 8),
    to_signed(3, 8),
    to_signed(2, 8),
    to_signed(1, 8),
    to_signed(0, 8),
    to_signed(0, 8),
    to_signed(-1, 8),
    to_signed(-2, 8),
    to_signed(-3, 8),
    to_signed(-4, 8),
    to_signed(-5, 8),
    to_signed(-6, 8),
    to_signed(-7, 8),
    to_signed(-6, 8),
    to_signed(-6, 8),
    to_signed(-6, 8),
    to_signed(-6, 8),
    to_signed(-5, 8),
    to_signed(-4, 8),
    to_signed(-4, 8),
    to_signed(-5, 8),
    to_signed(-7, 8),
    to_signed(-6, 8),
    to_signed(-5, 8),
    to_signed(-4, 8),
    to_signed(-4, 8),
    to_signed(-4, 8),
    to_signed(-5, 8),
    to_signed(-4, 8),
    to_signed(-4, 8),
    to_signed(-4, 8),
    to_signed(-3, 8),
    to_signed(-3, 8),
    to_signed(-3, 8),
    to_signed(-1, 8),
    to_signed(1, 8),
    to_signed(2, 8),
    to_signed(4, 8),
    to_signed(5, 8),
    to_signed(6, 8),
    to_signed(6, 8),
    to_signed(6, 8),
    to_signed(4, 8),
    to_signed(3, 8),
    to_signed(3, 8),
    to_signed(4, 8),
    to_signed(7, 8),
    to_signed(8, 8),
    to_signed(7, 8),
    to_signed(6, 8),
    to_signed(5, 8),
    to_signed(5, 8),
    to_signed(4, 8),
    to_signed(2, 8),
    to_signed(1, 8),
    to_signed(1, 8),
    to_signed(2, 8),
    to_signed(3, 8),
    to_signed(4, 8),
    to_signed(2, 8),
    to_signed(1, 8),
    to_signed(0, 8),
    to_signed(-1, 8),
    to_signed(-2, 8),
    to_signed(-4, 8),
    to_signed(-3, 8),
    to_signed(-2, 8),
    to_signed(-1, 8),
    to_signed(-2, 8),
    to_signed(-4, 8),
    to_signed(-4, 8),
    to_signed(-4, 8),
    to_signed(-4, 8),
    to_signed(-5, 8),
    to_signed(-5, 8),
    to_signed(-4, 8),
    to_signed(-4, 8),
    to_signed(-5, 8),
    to_signed(-6, 8),
    to_signed(-6, 8),
    to_signed(-5, 8),
    to_signed(-3, 8),
    to_signed(-3, 8),
    to_signed(-4, 8),
    to_signed(-5, 8),
    to_signed(-5, 8),
    to_signed(-5, 8),
    to_signed(-4, 8),
    to_signed(-3, 8),
    to_signed(-2, 8),
    to_signed(-2, 8),
    to_signed(-3, 8),
    to_signed(-2, 8),
    to_signed(-1, 8),
    to_signed(0, 8),
    to_signed(1, 8),
    to_signed(1, 8),
    to_signed(2, 8),
    to_signed(2, 8),
    to_signed(2, 8),
    to_signed(1, 8),
    to_signed(1, 8),
    to_signed(3, 8),
    to_signed(5, 8),
    to_signed(5, 8),
    to_signed(3, 8),
    to_signed(1, 8),
    to_signed(2, 8),
    to_signed(4, 8),
    to_signed(4, 8),
    to_signed(3, 8),
    to_signed(1, 8),
    to_signed(1, 8),
    to_signed(1, 8),
    to_signed(2, 8),
    to_signed(3, 8),
    to_signed(4, 8),
    to_signed(2, 8),
    to_signed(-2, 8),
    to_signed(-7, 8),
    to_signed(-9, 8),
    to_signed(-8, 8),
    to_signed(-6, 8),
    to_signed(-6, 8),
    to_signed(-5, 8),
    to_signed(-2, 8),
    to_signed(-1, 8),
    to_signed(-3, 8),
    to_signed(-6, 8),
    to_signed(-6, 8),
    to_signed(-4, 8),
    to_signed(-3, 8),
    to_signed(-5, 8),
    to_signed(-6, 8),
    to_signed(-6, 8),
    to_signed(-4, 8),
    to_signed(-4, 8),
    to_signed(-5, 8),
    to_signed(-8, 8),
    to_signed(-9, 8),
    to_signed(-9, 8),
    to_signed(-9, 8),
    to_signed(-9, 8),
    to_signed(-10, 8),
    to_signed(-9, 8),
    to_signed(-6, 8),
    to_signed(-3, 8),
    to_signed(-2, 8),
    to_signed(-5, 8),
    to_signed(-8, 8),
    to_signed(-8, 8),
    to_signed(-5, 8),
    to_signed(-2, 8),
    to_signed(-2, 8),
    to_signed(-4, 8),
    to_signed(-5, 8),
    to_signed(-3, 8),
    to_signed(-2, 8),
    to_signed(-2, 8),
    to_signed(-2, 8),
    to_signed(-2, 8),
    to_signed(-2, 8),
    to_signed(-2, 8),
    to_signed(-3, 8),
    to_signed(-5, 8),
    to_signed(-6, 8),
    to_signed(-6, 8),
    to_signed(-4, 8),
    to_signed(-1, 8),
    to_signed(-1, 8),
    to_signed(-3, 8),
    to_signed(-4, 8),
    to_signed(-4, 8),
    to_signed(-1, 8),
    to_signed(0, 8),
    to_signed(1, 8),
    to_signed(1, 8),
    to_signed(2, 8),
    to_signed(2, 8),
    to_signed(1, 8),
    to_signed(1, 8),
    to_signed(1, 8),
    to_signed(3, 8),
    to_signed(3, 8),
    to_signed(2, 8),
    to_signed(1, 8),
    to_signed(1, 8),
    to_signed(3, 8),
    to_signed(3, 8),
    to_signed(3, 8),
    to_signed(3, 8),
    to_signed(3, 8),
    to_signed(5, 8),
    to_signed(5, 8),
    to_signed(5, 8),
    to_signed(4, 8),
    to_signed(4, 8),
    to_signed(5, 8),
    to_signed(4, 8),
    to_signed(1, 8),
    to_signed(-1, 8),
    to_signed(-2, 8),
    to_signed(0, 8),
    to_signed(1, 8),
    to_signed(1, 8),
    to_signed(1, 8),
    to_signed(1, 8),
    to_signed(1, 8),
    to_signed(1, 8),
    to_signed(1, 8),
    to_signed(2, 8),
    to_signed(2, 8),
    to_signed(2, 8),
    to_signed(2, 8),
    to_signed(4, 8),
    to_signed(6, 8),
    to_signed(8, 8),
    to_signed(7, 8),
    to_signed(7, 8),
    to_signed(8, 8),
    to_signed(8, 8),
    to_signed(8, 8),
    to_signed(8, 8),
    to_signed(8, 8),
    to_signed(8, 8),
    to_signed(9, 8),
    to_signed(11, 8),
    to_signed(11, 8),
    to_signed(10, 8),
    to_signed(9, 8),
    to_signed(9, 8),
    to_signed(10, 8),
    to_signed(12, 8),
    to_signed(13, 8),
    to_signed(13, 8),
    to_signed(14, 8),
    to_signed(14, 8),
    to_signed(14, 8),
    to_signed(13, 8),
    to_signed(12, 8),
    to_signed(12, 8),
    to_signed(14, 8),
    to_signed(15, 8),
    to_signed(14, 8),
    to_signed(12, 8),
    to_signed(10, 8),
    to_signed(8, 8),
    to_signed(8, 8),
    to_signed(8, 8),
    to_signed(7, 8),
    to_signed(6, 8),
    to_signed(6, 8),
    to_signed(5, 8),
    to_signed(4, 8),
    to_signed(2, 8),
    to_signed(0, 8),
    to_signed(0, 8),
    to_signed(1, 8),
    to_signed(3, 8),
    to_signed(2, 8),
    to_signed(0, 8),
    to_signed(-1, 8),
    to_signed(-1, 8),
    to_signed(-3, 8),
    to_signed(-4, 8),
    to_signed(-5, 8),
    to_signed(-6, 8),
    to_signed(-7, 8),
    to_signed(-8, 8),
    to_signed(-9, 8),
    to_signed(-8, 8),
    to_signed(-8, 8),
    to_signed(-6, 8),
    to_signed(-6, 8),
    to_signed(-8, 8),
    to_signed(-10, 8),
    to_signed(-10, 8),
    to_signed(-9, 8),
    to_signed(-8, 8),
    to_signed(-8, 8),
    to_signed(-6, 8),
    to_signed(-3, 8),
    to_signed(-1, 8),
    to_signed(-1, 8),
    to_signed(-2, 8),
    to_signed(-3, 8),
    to_signed(-2, 8),
    to_signed(-2, 8),
    to_signed(-2, 8),
    to_signed(-2, 8),
    to_signed(-1, 8),
    to_signed(3, 8),
    to_signed(5, 8),
    to_signed(5, 8),
    to_signed(5, 8),
    to_signed(4, 8),
    to_signed(5, 8),
    to_signed(5, 8),
    to_signed(5, 8),
    to_signed(5, 8),
    to_signed(4, 8),
    to_signed(3, 8),
    to_signed(2, 8),
    to_signed(1, 8),
    to_signed(1, 8),
    to_signed(1, 8),
    to_signed(0, 8),
    to_signed(-1, 8),
    to_signed(-1, 8),
    to_signed(-1, 8),
    to_signed(-3, 8),
    to_signed(-4, 8),
    to_signed(-4, 8),
    to_signed(-5, 8),
    to_signed(-6, 8),
    to_signed(-8, 8),
    to_signed(-10, 8),
    to_signed(-11, 8),
    to_signed(-12, 8),
    to_signed(-12, 8),
    to_signed(-12, 8),
    to_signed(-12, 8),
    to_signed(-12, 8),
    to_signed(-12, 8),
    to_signed(-12, 8),
    to_signed(-11, 8),
    to_signed(-10, 8),
    to_signed(-10, 8),
    to_signed(-11, 8),
    to_signed(-12, 8),
    to_signed(-12, 8),
    to_signed(-12, 8),
    to_signed(-11, 8),
    to_signed(-11, 8),
    to_signed(-12, 8),
    to_signed(-13, 8),
    to_signed(-12, 8),
    to_signed(-9, 8),
    to_signed(-7, 8),
    to_signed(-7, 8),
    to_signed(-6, 8),
    to_signed(-4, 8),
    to_signed(-3, 8),
    to_signed(-4, 8),
    to_signed(-5, 8),
    to_signed(-4, 8),
    to_signed(-2, 8),
    to_signed(0, 8),
    to_signed(0, 8),
    to_signed(1, 8),
    to_signed(2, 8),
    to_signed(4, 8),
    to_signed(6, 8),
    to_signed(6, 8),
    to_signed(6, 8),
    to_signed(5, 8),
    to_signed(5, 8),
    to_signed(4, 8),
    to_signed(4, 8),
    to_signed(5, 8),
    to_signed(6, 8),
    to_signed(7, 8),
    to_signed(6, 8),
    to_signed(6, 8),
    to_signed(4, 8),
    to_signed(2, 8),
    to_signed(1, 8),
    to_signed(2, 8),
    to_signed(2, 8),
    to_signed(3, 8),
    to_signed(3, 8),
    to_signed(4, 8),
    to_signed(3, 8),
    to_signed(2, 8),
    to_signed(0, 8),
    to_signed(-1, 8),
    to_signed(-3, 8),
    to_signed(-3, 8),
    to_signed(-4, 8),
    to_signed(-4, 8),
    to_signed(-4, 8),
    to_signed(-5, 8),
    to_signed(-5, 8),
    to_signed(-6, 8),
    to_signed(-6, 8),
    to_signed(-6, 8),
    to_signed(-7, 8),
    to_signed(-7, 8),
    to_signed(-6, 8),
    to_signed(-6, 8),
    to_signed(-6, 8),
    to_signed(-6, 8),
    to_signed(-5, 8),
    to_signed(-4, 8),
    to_signed(-3, 8),
    to_signed(-2, 8),
    to_signed(-2, 8),
    to_signed(-3, 8),
    to_signed(-3, 8),
    to_signed(-2, 8),
    to_signed(-2, 8),
    to_signed(-3, 8),
    to_signed(-2, 8),
    to_signed(0, 8),
    to_signed(2, 8),
    to_signed(3, 8),
    to_signed(4, 8),
    to_signed(5, 8),
    to_signed(7, 8),
    to_signed(8, 8),
    to_signed(8, 8),
    to_signed(8, 8),
    to_signed(9, 8),
    to_signed(11, 8),
    to_signed(12, 8),
    to_signed(13, 8),
    to_signed(13, 8),
    to_signed(15, 8),
    to_signed(16, 8),
    to_signed(15, 8),
    to_signed(13, 8),
    to_signed(12, 8),
    to_signed(12, 8),
    to_signed(14, 8),
    to_signed(14, 8),
    to_signed(14, 8),
    to_signed(14, 8),
    to_signed(13, 8),
    to_signed(13, 8),
    to_signed(13, 8),
    to_signed(12, 8),
    to_signed(12, 8),
    to_signed(10, 8),
    to_signed(9, 8),
    to_signed(9, 8),
    to_signed(9, 8),
    to_signed(8, 8),
    to_signed(8, 8),
    to_signed(7, 8),
    to_signed(6, 8),
    to_signed(4, 8),
    to_signed(2, 8),
    to_signed(1, 8),
    to_signed(0, 8),
    to_signed(-1, 8),
    to_signed(0, 8),
    to_signed(0, 8),
    to_signed(0, 8),
    to_signed(1, 8),
    to_signed(1, 8),
    to_signed(0, 8),
    to_signed(-2, 8),
    to_signed(-3, 8),
    to_signed(-3, 8),
    to_signed(-2, 8),
    to_signed(-1, 8),
    to_signed(0, 8),
    to_signed(1, 8),
    to_signed(1, 8),
    to_signed(0, 8),
    to_signed(1, 8),
    to_signed(2, 8),
    to_signed(2, 8),
    to_signed(2, 8),
    to_signed(2, 8),
    to_signed(2, 8),
    to_signed(2, 8),
    to_signed(2, 8),
    to_signed(2, 8),
    to_signed(3, 8),
    to_signed(4, 8),
    to_signed(4, 8),
    to_signed(4, 8),
    to_signed(4, 8),
    to_signed(3, 8),
    to_signed(4, 8),
    to_signed(4, 8),
    to_signed(5, 8),
    to_signed(6, 8),
    to_signed(5, 8),
    to_signed(4, 8),
    to_signed(3, 8),
    to_signed(3, 8),
    to_signed(3, 8),
    to_signed(2, 8),
    to_signed(1, 8),
    to_signed(-1, 8),
    to_signed(-3, 8),
    to_signed(-4, 8),
    to_signed(-6, 8),
    to_signed(-7, 8),
    to_signed(-7, 8),
    to_signed(-8, 8),
    to_signed(-8, 8),
    to_signed(-8, 8),
    to_signed(-8, 8),
    to_signed(-8, 8),
    to_signed(-10, 8),
    to_signed(-12, 8),
    to_signed(-13, 8),
    to_signed(-13, 8),
    to_signed(-13, 8),
    to_signed(-12, 8),
    to_signed(-12, 8),
    to_signed(-13, 8),
    to_signed(-14, 8),
    to_signed(-14, 8),
    to_signed(-15, 8),
    to_signed(-16, 8),
    to_signed(-17, 8),
    to_signed(-17, 8),
    to_signed(-17, 8),
    to_signed(-17, 8),
    to_signed(-18, 8),
    to_signed(-17, 8),
    to_signed(-15, 8),
    to_signed(-14, 8),
    to_signed(-15, 8),
    to_signed(-16, 8),
    to_signed(-16, 8),
    to_signed(-14, 8),
    to_signed(-12, 8),
    to_signed(-11, 8),
    to_signed(-9, 8),
    to_signed(-8, 8),
    to_signed(-7, 8),
    to_signed(-7, 8),
    to_signed(-9, 8),
    to_signed(-9, 8),
    to_signed(-8, 8),
    to_signed(-6, 8),
    to_signed(-4, 8),
    to_signed(-3, 8),
    to_signed(-2, 8),
    to_signed(-2, 8),
    to_signed(-2, 8),
    to_signed(-2, 8),
    to_signed(-1, 8),
    to_signed(0, 8),
    to_signed(1, 8),
    to_signed(3, 8),
    to_signed(4, 8),
    to_signed(4, 8),
    to_signed(4, 8),
    to_signed(5, 8),
    to_signed(5, 8),
    to_signed(5, 8),
    to_signed(4, 8),
    to_signed(3, 8),
    to_signed(2, 8),
    to_signed(1, 8),
    to_signed(0, 8),
    to_signed(-2, 8),
    to_signed(-3, 8),
    to_signed(-3, 8),
    to_signed(-3, 8),
    to_signed(-3, 8),
    to_signed(-4, 8),
    to_signed(-6, 8),
    to_signed(-7, 8),
    to_signed(-6, 8),
    to_signed(-6, 8),
    to_signed(-7, 8),
    to_signed(-9, 8),
    to_signed(-9, 8),
    to_signed(-7, 8),
    to_signed(-6, 8),
    to_signed(-6, 8),
    to_signed(-7, 8),
    to_signed(-7, 8),
    to_signed(-6, 8),
    to_signed(-6, 8),
    to_signed(-8, 8),
    to_signed(-9, 8),
    to_signed(-10, 8),
    to_signed(-8, 8),
    to_signed(-7, 8),
    to_signed(-7, 8),
    to_signed(-7, 8),
    to_signed(-5, 8),
    to_signed(-3, 8),
    to_signed(-1, 8),
    to_signed(1, 8),
    to_signed(1, 8),
    to_signed(2, 8),
    to_signed(2, 8),
    to_signed(3, 8),
    to_signed(4, 8),
    to_signed(4, 8),
    to_signed(4, 8),
    to_signed(4, 8),
    to_signed(4, 8),
    to_signed(5, 8),
    to_signed(5, 8),
    to_signed(4, 8),
    to_signed(4, 8),
    to_signed(4, 8),
    to_signed(5, 8),
    to_signed(6, 8),
    to_signed(7, 8),
    to_signed(6, 8),
    to_signed(5, 8),
    to_signed(6, 8),
    to_signed(7, 8),
    to_signed(7, 8),
    to_signed(7, 8),
    to_signed(7, 8),
    to_signed(6, 8),
    to_signed(6, 8),
    to_signed(5, 8),
    to_signed(5, 8),
    to_signed(5, 8),
    to_signed(4, 8),
    to_signed(3, 8),
    to_signed(2, 8),
    to_signed(0, 8),
    to_signed(-2, 8),
    to_signed(-3, 8),
    to_signed(-4, 8),
    to_signed(-5, 8),
    to_signed(-6, 8),
    to_signed(-6, 8),
    to_signed(-6, 8),
    to_signed(-6, 8),
    to_signed(-7, 8),
    to_signed(-7, 8),
    to_signed(-6, 8),
    to_signed(-5, 8),
    to_signed(-5, 8),
    to_signed(-5, 8),
    to_signed(-3, 8),
    to_signed(-2, 8),
    to_signed(-1, 8),
    to_signed(-1, 8),
    to_signed(-1, 8),
    to_signed(-2, 8),
    to_signed(-3, 8),
    to_signed(-2, 8),
    to_signed(-1, 8),
    to_signed(0, 8),
    to_signed(1, 8),
    to_signed(1, 8),
    to_signed(1, 8),
    to_signed(2, 8),
    to_signed(3, 8),
    to_signed(3, 8),
    to_signed(3, 8),
    to_signed(3, 8),
    to_signed(4, 8),
    to_signed(5, 8),
    to_signed(6, 8),
    to_signed(8, 8),
    to_signed(9, 8),
    to_signed(10, 8),
    to_signed(8, 8),
    to_signed(6, 8),
    to_signed(4, 8),
    to_signed(3, 8),
    to_signed(3, 8),
    to_signed(3, 8),
    to_signed(3, 8),
    to_signed(2, 8),
    to_signed(1, 8),
    to_signed(-1, 8),
    to_signed(-2, 8),
    to_signed(-2, 8),
    to_signed(0, 8),
    to_signed(1, 8),
    to_signed(1, 8),
    to_signed(0, 8),
    to_signed(-1, 8),
    to_signed(0, 8),
    to_signed(0, 8),
    to_signed(0, 8),
    to_signed(-1, 8),
    to_signed(-1, 8),
    to_signed(-2, 8),
    to_signed(-2, 8),
    to_signed(-3, 8),
    to_signed(-4, 8),
    to_signed(-4, 8),
    to_signed(-3, 8),
    to_signed(-2, 8),
    to_signed(-3, 8),
    to_signed(-5, 8),
    to_signed(-7, 8),
    to_signed(-7, 8),
    to_signed(-6, 8),
    to_signed(-6, 8),
    to_signed(-7, 8),
    to_signed(-7, 8),
    to_signed(-6, 8),
    to_signed(-5, 8),
    to_signed(-3, 8),
    to_signed(-3, 8),
    to_signed(-4, 8),
    to_signed(-6, 8),
    to_signed(-6, 8),
    to_signed(-5, 8),
    to_signed(-4, 8),
    to_signed(-5, 8),
    to_signed(-7, 8),
    to_signed(-8, 8),
    to_signed(-8, 8),
    to_signed(-7, 8),
    to_signed(-6, 8),
    to_signed(-5, 8),
    to_signed(-5, 8),
    to_signed(-4, 8),
    to_signed(-3, 8),
    to_signed(-3, 8),
    to_signed(-5, 8),
    to_signed(-5, 8),
    to_signed(-3, 8),
    to_signed(-1, 8),
    to_signed(-1, 8),
    to_signed(0, 8),
    to_signed(1, 8),
    to_signed(3, 8),
    to_signed(2, 8),
    to_signed(1, 8),
    to_signed(0, 8),
    to_signed(1, 8),
    to_signed(1, 8),
    to_signed(1, 8),
    to_signed(0, 8),
    to_signed(-2, 8),
    to_signed(-3, 8),
    to_signed(-4, 8),
    to_signed(-5, 8),
    to_signed(-6, 8),
    to_signed(-6, 8),
    to_signed(-5, 8),
    to_signed(-3, 8),
    to_signed(-3, 8),
    to_signed(-3, 8),
    to_signed(-2, 8),
    to_signed(-2, 8),
    to_signed(-2, 8),
    to_signed(-2, 8),
    to_signed(-2, 8),
    to_signed(-2, 8),
    to_signed(-3, 8),
    to_signed(-4, 8),
    to_signed(-5, 8),
    to_signed(-5, 8),
    to_signed(-4, 8),
    to_signed(-2, 8),
    to_signed(0, 8),
    to_signed(0, 8),
    to_signed(0, 8),
    to_signed(0, 8),
    to_signed(1, 8),
    to_signed(3, 8),
    to_signed(5, 8),
    to_signed(7, 8),
    to_signed(7, 8),
    to_signed(7, 8),
    to_signed(8, 8),
    to_signed(11, 8),
    to_signed(14, 8),
    to_signed(15, 8),
    to_signed(16, 8),
    to_signed(16, 8),
    to_signed(15, 8),
    to_signed(16, 8),
    to_signed(18, 8),
    to_signed(20, 8),
    to_signed(22, 8),
    to_signed(21, 8),
    to_signed(20, 8),
    to_signed(18, 8),
    to_signed(17, 8),
    to_signed(16, 8),
    to_signed(16, 8),
    to_signed(16, 8),
    to_signed(16, 8),
    to_signed(16, 8),
    to_signed(15, 8),
    to_signed(15, 8),
    to_signed(15, 8),
    to_signed(15, 8),
    to_signed(15, 8),
    to_signed(15, 8),
    to_signed(13, 8),
    to_signed(11, 8),
    to_signed(9, 8),
    to_signed(7, 8),
    to_signed(6, 8),
    to_signed(6, 8),
    to_signed(5, 8),
    to_signed(4, 8),
    to_signed(2, 8),
    to_signed(1, 8),
    to_signed(-1, 8),
    to_signed(-2, 8),
    to_signed(-3, 8),
    to_signed(-3, 8),
    to_signed(-4, 8),
    to_signed(-7, 8),
    to_signed(-8, 8),
    to_signed(-7, 8),
    to_signed(-6, 8),
    to_signed(-4, 8),
    to_signed(-3, 8),
    to_signed(-3, 8),
    to_signed(-4, 8),
    to_signed(-4, 8),
    to_signed(-4, 8),
    to_signed(-4, 8),
    to_signed(-4, 8),
    to_signed(-4, 8),
    to_signed(-3, 8),
    to_signed(-3, 8),
    to_signed(-3, 8),
    to_signed(-3, 8),
    to_signed(-3, 8),
    to_signed(-3, 8),
    to_signed(-3, 8),
    to_signed(-2, 8),
    to_signed(0, 8),
    to_signed(2, 8),
    to_signed(4, 8),
    to_signed(4, 8),
    to_signed(5, 8),
    to_signed(6, 8),
    to_signed(6, 8),
    to_signed(7, 8),
    to_signed(8, 8),
    to_signed(9, 8),
    to_signed(8, 8),
    to_signed(7, 8),
    to_signed(6, 8),
    to_signed(6, 8),
    to_signed(6, 8),
    to_signed(6, 8),
    to_signed(7, 8),
    to_signed(6, 8),
    to_signed(5, 8),
    to_signed(3, 8),
    to_signed(3, 8),
    to_signed(3, 8),
    to_signed(4, 8),
    to_signed(4, 8),
    to_signed(5, 8),
    to_signed(5, 8),
    to_signed(6, 8),
    to_signed(6, 8),
    to_signed(5, 8),
    to_signed(4, 8),
    to_signed(3, 8),
    to_signed(3, 8),
    to_signed(2, 8),
    to_signed(0, 8),
    to_signed(-1, 8),
    to_signed(-1, 8),
    to_signed(-1, 8),
    to_signed(-2, 8),
    to_signed(-3, 8),
    to_signed(-4, 8),
    to_signed(-5, 8),
    to_signed(-5, 8),
    to_signed(-6, 8),
    to_signed(-7, 8),
    to_signed(-6, 8),
    to_signed(-5, 8),
    to_signed(-3, 8),
    to_signed(-3, 8),
    to_signed(-4, 8),
    to_signed(-4, 8),
    to_signed(-3, 8),
    to_signed(-3, 8),
    to_signed(-3, 8),
    to_signed(-3, 8),
    to_signed(-2, 8),
    to_signed(-2, 8),
    to_signed(-2, 8),
    to_signed(-1, 8),
    to_signed(0, 8),
    to_signed(-1, 8),
    to_signed(-2, 8),
    to_signed(-3, 8),
    to_signed(-3, 8),
    to_signed(-3, 8),
    to_signed(-3, 8),
    to_signed(-3, 8),
    to_signed(-3, 8),
    to_signed(-2, 8),
    to_signed(-2, 8),
    to_signed(-2, 8),
    to_signed(-2, 8),
    to_signed(-2, 8),
    to_signed(0, 8),
    to_signed(-1, 8),
    to_signed(-2, 8),
    to_signed(-3, 8),
    to_signed(-3, 8),
    to_signed(-3, 8),
    to_signed(-4, 8),
    to_signed(-5, 8),
    to_signed(-6, 8),
    to_signed(-8, 8),
    to_signed(-9, 8),
    to_signed(-11, 8),
    to_signed(-13, 8),
    to_signed(-13, 8),
    to_signed(-14, 8),
    to_signed(-15, 8),
    to_signed(-15, 8),
    to_signed(-16, 8),
    to_signed(-15, 8),
    to_signed(-13, 8),
    to_signed(-13, 8),
    to_signed(-13, 8),
    to_signed(-13, 8),
    to_signed(-12, 8),
    to_signed(-12, 8),
    to_signed(-12, 8),
    to_signed(-12, 8),
    to_signed(-12, 8),
    to_signed(-13, 8),
    to_signed(-15, 8),
    to_signed(-15, 8),
    to_signed(-14, 8),
    to_signed(-12, 8),
    to_signed(-13, 8),
    to_signed(-14, 8),
    to_signed(-13, 8),
    to_signed(-11, 8),
    to_signed(-10, 8),
    to_signed(-8, 8),
    to_signed(-7, 8),
    to_signed(-5, 8),
    to_signed(-4, 8),
    to_signed(-3, 8),
    to_signed(-3, 8),
    to_signed(-1, 8),
    to_signed(2, 8),
    to_signed(5, 8),
    to_signed(5, 8),
    to_signed(5, 8),
    to_signed(5, 8),
    to_signed(5, 8),
    to_signed(6, 8),
    to_signed(7, 8),
    to_signed(7, 8),
    to_signed(7, 8),
    to_signed(6, 8),
    to_signed(4, 8),
    to_signed(3, 8),
    to_signed(4, 8),
    to_signed(6, 8),
    to_signed(7, 8),
    to_signed(8, 8),
    to_signed(8, 8),
    to_signed(9, 8),
    to_signed(8, 8),
    to_signed(7, 8),
    to_signed(6, 8),
    to_signed(6, 8),
    to_signed(7, 8),
    to_signed(8, 8),
    to_signed(8, 8),
    to_signed(7, 8),
    to_signed(4, 8),
    to_signed(3, 8),
    to_signed(1, 8),
    to_signed(-1, 8),
    to_signed(-3, 8),
    to_signed(-3, 8),
    to_signed(-3, 8),
    to_signed(-4, 8),
    to_signed(-4, 8),
    to_signed(-4, 8),
    to_signed(-4, 8),
    to_signed(-4, 8),
    to_signed(-5, 8),
    to_signed(-5, 8),
    to_signed(-5, 8),
    to_signed(-5, 8),
    to_signed(-6, 8),
    to_signed(-6, 8),
    to_signed(-6, 8),
    to_signed(-6, 8),
    to_signed(-6, 8),
    to_signed(-7, 8),
    to_signed(-8, 8),
    to_signed(-8, 8),
    to_signed(-8, 8),
    to_signed(-8, 8),
    to_signed(-8, 8),
    to_signed(-9, 8),
    to_signed(-10, 8),
    to_signed(-9, 8),
    to_signed(-8, 8),
    to_signed(-7, 8),
    to_signed(-6, 8),
    to_signed(-4, 8),
    to_signed(-3, 8),
    to_signed(-2, 8),
    to_signed(-2, 8),
    to_signed(-1, 8),
    to_signed(1, 8),
    to_signed(3, 8),
    to_signed(4, 8),
    to_signed(4, 8),
    to_signed(3, 8),
    to_signed(2, 8),
    to_signed(1, 8),
    to_signed(0, 8),
    to_signed(-1, 8),
    to_signed(-1, 8),
    to_signed(-1, 8),
    to_signed(-1, 8),
    to_signed(-2, 8),
    to_signed(-4, 8),
    to_signed(-5, 8),
    to_signed(-6, 8),
    to_signed(-5, 8),
    to_signed(-5, 8),
    to_signed(-5, 8),
    to_signed(-6, 8),
    to_signed(-6, 8),
    to_signed(-6, 8),
    to_signed(-5, 8),
    to_signed(-6, 8),
    to_signed(-6, 8),
    to_signed(-7, 8),
    to_signed(-9, 8),
    to_signed(-10, 8),
    to_signed(-11, 8),
    to_signed(-11, 8),
    to_signed(-11, 8),
    to_signed(-11, 8),
    to_signed(-10, 8),
    to_signed(-11, 8),
    to_signed(-13, 8),
    to_signed(-15, 8),
    to_signed(-16, 8),
    to_signed(-14, 8),
    to_signed(-13, 8),
    to_signed(-13, 8),
    to_signed(-12, 8),
    to_signed(-10, 8),
    to_signed(-9, 8),
    to_signed(-9, 8),
    to_signed(-9, 8),
    to_signed(-8, 8),
    to_signed(-6, 8),
    to_signed(-5, 8),
    to_signed(-4, 8),
    to_signed(-5, 8),
    to_signed(-6, 8),
    to_signed(-7, 8),
    to_signed(-7, 8),
    to_signed(-7, 8),
    to_signed(-6, 8),
    to_signed(-4, 8),
    to_signed(-3, 8),
    to_signed(-3, 8),
    to_signed(-3, 8),
    to_signed(-1, 8),
    to_signed(1, 8),
    to_signed(4, 8),
    to_signed(7, 8),
    to_signed(9, 8),
    to_signed(10, 8),
    to_signed(10, 8),
    to_signed(10, 8),
    to_signed(10, 8),
    to_signed(10, 8),
    to_signed(10, 8),
    to_signed(11, 8),
    to_signed(13, 8),
    to_signed(14, 8),
    to_signed(15, 8),
    to_signed(14, 8),
    to_signed(14, 8),
    to_signed(13, 8),
    to_signed(13, 8),
    to_signed(14, 8),
    to_signed(14, 8),
    to_signed(13, 8),
    to_signed(11, 8),
    to_signed(9, 8),
    to_signed(9, 8),
    to_signed(8, 8),
    to_signed(8, 8),
    to_signed(8, 8),
    to_signed(8, 8),
    to_signed(9, 8),
    to_signed(9, 8),
    to_signed(10, 8),
    to_signed(9, 8),
    to_signed(8, 8),
    to_signed(6, 8),
    to_signed(4, 8),
    to_signed(4, 8),
    to_signed(4, 8),
    to_signed(5, 8),
    to_signed(4, 8),
    to_signed(3, 8),
    to_signed(0, 8),
    to_signed(-2, 8),
    to_signed(-3, 8),
    to_signed(-4, 8),
    to_signed(-4, 8),
    to_signed(-3, 8),
    to_signed(-2, 8),
    to_signed(-1, 8),
    to_signed(0, 8),
    to_signed(1, 8),
    to_signed(1, 8),
    to_signed(2, 8),
    to_signed(2, 8),
    to_signed(1, 8),
    to_signed(0, 8),
    to_signed(0, 8),
    to_signed(-1, 8),
    to_signed(-1, 8),
    to_signed(-1, 8),
    to_signed(-2, 8),
    to_signed(-3, 8),
    to_signed(-4, 8),
    to_signed(-5, 8),
    to_signed(-5, 8),
    to_signed(-5, 8),
    to_signed(-3, 8),
    to_signed(0, 8),
    to_signed(3, 8),
    to_signed(4, 8),
    to_signed(5, 8),
    to_signed(5, 8),
    to_signed(6, 8),
    to_signed(7, 8),
    to_signed(8, 8),
    to_signed(8, 8),
    to_signed(9, 8),
    to_signed(10, 8),
    to_signed(11, 8),
    to_signed(10, 8),
    to_signed(9, 8),
    to_signed(7, 8),
    to_signed(7, 8),
    to_signed(7, 8),
    to_signed(7, 8),
    to_signed(6, 8),
    to_signed(5, 8),
    to_signed(5, 8),
    to_signed(6, 8),
    to_signed(7, 8),
    to_signed(7, 8),
    to_signed(8, 8),
    to_signed(8, 8),
    to_signed(8, 8),
    to_signed(7, 8),
    to_signed(6, 8),
    to_signed(6, 8),
    to_signed(5, 8),
    to_signed(5, 8),
    to_signed(4, 8),
    to_signed(2, 8),
    to_signed(1, 8),
    to_signed(0, 8),
    to_signed(0, 8),
    to_signed(0, 8),
    to_signed(-1, 8),
    to_signed(-2, 8),
    to_signed(-5, 8),
    to_signed(-7, 8),
    to_signed(-9, 8),
    to_signed(-9, 8),
    to_signed(-7, 8),
    to_signed(-6, 8),
    to_signed(-5, 8),
    to_signed(-5, 8),
    to_signed(-5, 8),
    to_signed(-4, 8),
    to_signed(-4, 8),
    to_signed(-4, 8),
    to_signed(-3, 8),
    to_signed(-3, 8),
    to_signed(-3, 8),
    to_signed(-3, 8),
    to_signed(-4, 8),
    to_signed(-6, 8),
    to_signed(-8, 8),
    to_signed(-8, 8),
    to_signed(-8, 8),
    to_signed(-7, 8),
    to_signed(-6, 8),
    to_signed(-6, 8),
    to_signed(-6, 8),
    to_signed(-7, 8),
    to_signed(-6, 8),
    to_signed(-5, 8),
    to_signed(-4, 8),
    to_signed(-2, 8),
    to_signed(0, 8),
    to_signed(0, 8),
    to_signed(0, 8),
    to_signed(-1, 8),
    to_signed(0, 8),
    to_signed(0, 8),
    to_signed(0, 8),
    to_signed(0, 8),
    to_signed(0, 8),
    to_signed(0, 8),
    to_signed(-1, 8),
    to_signed(-1, 8),
    to_signed(-2, 8),
    to_signed(-2, 8),
    to_signed(-2, 8),
    to_signed(-1, 8),
    to_signed(-1, 8),
    to_signed(-1, 8),
    to_signed(0, 8),
    to_signed(2, 8),
    to_signed(3, 8),
    to_signed(4, 8),
    to_signed(3, 8),
    to_signed(2, 8),
    to_signed(2, 8),
    to_signed(3, 8),
    to_signed(3, 8),
    to_signed(3, 8),
    to_signed(3, 8),
    to_signed(2, 8),
    to_signed(2, 8),
    to_signed(1, 8),
    to_signed(1, 8),
    to_signed(0, 8),
    to_signed(-1, 8),
    to_signed(-2, 8),
    to_signed(-3, 8),
    to_signed(-3, 8),
    to_signed(-3, 8),
    to_signed(-2, 8),
    to_signed(-1, 8),
    to_signed(1, 8),
    to_signed(1, 8),
    to_signed(1, 8),
    to_signed(1, 8),
    to_signed(0, 8),
    to_signed(0, 8),
    to_signed(1, 8),
    to_signed(2, 8),
    to_signed(3, 8),
    to_signed(3, 8),
    to_signed(3, 8),
    to_signed(2, 8),
    to_signed(1, 8),
    to_signed(1, 8),
    to_signed(0, 8),
    to_signed(-1, 8),
    to_signed(-1, 8),
    to_signed(-1, 8),
    to_signed(-1, 8),
    to_signed(-2, 8),
    to_signed(-2, 8),
    to_signed(-1, 8),
    to_signed(-1, 8),
    to_signed(1, 8),
    to_signed(2, 8),
    to_signed(3, 8),
    to_signed(4, 8),
    to_signed(4, 8),
    to_signed(4, 8),
    to_signed(3, 8),
    to_signed(2, 8),
    to_signed(1, 8),
    to_signed(1, 8),
    to_signed(0, 8),
    to_signed(-1, 8),
    to_signed(-2, 8),
    to_signed(-3, 8),
    to_signed(-4, 8),
    to_signed(-5, 8),
    to_signed(-7, 8),
    to_signed(-8, 8),
    to_signed(-9, 8),
    to_signed(-8, 8),
    to_signed(-8, 8),
    to_signed(-7, 8),
    to_signed(-7, 8),
    to_signed(-7, 8),
    to_signed(-6, 8),
    to_signed(-6, 8),
    to_signed(-6, 8),
    to_signed(-7, 8),
    to_signed(-7, 8),
    to_signed(-7, 8),
    to_signed(-7, 8),
    to_signed(-8, 8),
    to_signed(-8, 8),
    to_signed(-9, 8),
    to_signed(-9, 8),
    to_signed(-10, 8),
    to_signed(-11, 8),
    to_signed(-12, 8),
    to_signed(-10, 8),
    to_signed(-8, 8),
    to_signed(-8, 8),
    to_signed(-9, 8),
    to_signed(-9, 8),
    to_signed(-8, 8),
    to_signed(-7, 8),
    to_signed(-6, 8),
    to_signed(-5, 8),
    to_signed(-4, 8),
    to_signed(-3, 8),
    to_signed(-3, 8),
    to_signed(-3, 8),
    to_signed(-2, 8),
    to_signed(-2, 8),
    to_signed(-2, 8),
    to_signed(-2, 8),
    to_signed(-2, 8),
    to_signed(-2, 8),
    to_signed(-1, 8),
    to_signed(-1, 8),
    to_signed(-1, 8),
    to_signed(-1, 8),
    to_signed(-1, 8),
    to_signed(-2, 8),
    to_signed(-2, 8),
    to_signed(-1, 8),
    to_signed(1, 8),
    to_signed(2, 8),
    to_signed(4, 8),
    to_signed(6, 8),
    to_signed(6, 8),
    to_signed(4, 8),
    to_signed(3, 8),
    to_signed(3, 8),
    to_signed(4, 8),
    to_signed(4, 8),
    to_signed(4, 8),
    to_signed(2, 8),
    to_signed(1, 8),
    to_signed(0, 8),
    to_signed(-1, 8),
    to_signed(-2, 8),
    to_signed(-2, 8),
    to_signed(-1, 8),
    to_signed(0, 8),
    to_signed(-1, 8),
    to_signed(-1, 8),
    to_signed(-2, 8),
    to_signed(-2, 8),
    to_signed(-2, 8),
    to_signed(-2, 8),
    to_signed(-2, 8),
    to_signed(-1, 8),
    to_signed(-1, 8),
    to_signed(0, 8),
    to_signed(0, 8),
    to_signed(-1, 8),
    to_signed(-2, 8),
    to_signed(-3, 8),
    to_signed(-4, 8),
    to_signed(-5, 8),
    to_signed(-5, 8),
    to_signed(-6, 8),
    to_signed(-5, 8),
    to_signed(-6, 8),
    to_signed(-7, 8),
    to_signed(-8, 8),
    to_signed(-9, 8),
    to_signed(-9, 8),
    to_signed(-9, 8),
    to_signed(-9, 8),
    to_signed(-8, 8),
    to_signed(-6, 8),
    to_signed(-4, 8),
    to_signed(-3, 8),
    to_signed(-2, 8),
    to_signed(-2, 8),
    to_signed(-2, 8),
    to_signed(-3, 8),
    to_signed(-3, 8),
    to_signed(-2, 8),
    to_signed(-2, 8),
    to_signed(-3, 8),
    to_signed(-4, 8),
    to_signed(-5, 8),
    to_signed(-6, 8),
    to_signed(-6, 8),
    to_signed(-5, 8),
    to_signed(-3, 8),
    to_signed(0, 8),
    to_signed(2, 8),
    to_signed(2, 8),
    to_signed(2, 8),
    to_signed(2, 8),
    to_signed(3, 8),
    to_signed(4, 8),
    to_signed(6, 8),
    to_signed(7, 8),
    to_signed(9, 8),
    to_signed(10, 8),
    to_signed(10, 8),
    to_signed(9, 8),
    to_signed(8, 8),
    to_signed(7, 8),
    to_signed(7, 8),
    to_signed(7, 8),
    to_signed(7, 8),
    to_signed(7, 8),
    to_signed(7, 8),
    to_signed(8, 8),
    to_signed(8, 8),
    to_signed(7, 8),
    to_signed(6, 8),
    to_signed(5, 8),
    to_signed(5, 8),
    to_signed(5, 8),
    to_signed(4, 8),
    to_signed(5, 8),
    to_signed(5, 8),
    to_signed(6, 8),
    to_signed(6, 8),
    to_signed(5, 8),
    to_signed(5, 8),
    to_signed(5, 8),
    to_signed(4, 8),
    to_signed(2, 8),
    to_signed(1, 8),
    to_signed(0, 8),
    to_signed(-1, 8),
    to_signed(-2, 8),
    to_signed(-4, 8),
    to_signed(-5, 8),
    to_signed(-5, 8),
    to_signed(-4, 8),
    to_signed(-4, 8),
    to_signed(-4, 8),
    to_signed(-4, 8),
    to_signed(-4, 8),
    to_signed(-4, 8),
    to_signed(-3, 8),
    to_signed(-3, 8),
    to_signed(-2, 8),
    to_signed(-1, 8),
    to_signed(-1, 8),
    to_signed(0, 8),
    to_signed(0, 8),
    to_signed(-1, 8),
    to_signed(-2, 8),
    to_signed(-3, 8),
    to_signed(-3, 8),
    to_signed(-4, 8),
    to_signed(-3, 8),
    to_signed(-2, 8),
    to_signed(-1, 8),
    to_signed(0, 8),
    to_signed(0, 8),
    to_signed(0, 8),
    to_signed(1, 8),
    to_signed(2, 8),
    to_signed(3, 8),
    to_signed(4, 8),
    to_signed(5, 8),
    to_signed(7, 8),
    to_signed(8, 8),
    to_signed(10, 8),
    to_signed(10, 8),
    to_signed(10, 8),
    to_signed(10, 8),
    to_signed(9, 8),
    to_signed(9, 8),
    to_signed(9, 8),
    to_signed(8, 8),
    to_signed(7, 8),
    to_signed(6, 8),
    to_signed(5, 8),
    to_signed(6, 8),
    to_signed(7, 8),
    to_signed(7, 8),
    to_signed(7, 8),
    to_signed(6, 8),
    to_signed(5, 8),
    to_signed(4, 8),
    to_signed(4, 8),
    to_signed(5, 8),
    to_signed(6, 8),
    to_signed(7, 8),
    to_signed(7, 8),
    to_signed(7, 8),
    to_signed(6, 8),
    to_signed(4, 8),
    to_signed(1, 8),
    to_signed(-1, 8),
    to_signed(-3, 8),
    to_signed(-4, 8),
    to_signed(-4, 8),
    to_signed(-5, 8),
    to_signed(-6, 8),
    to_signed(-7, 8),
    to_signed(-6, 8),
    to_signed(-6, 8),
    to_signed(-5, 8),
    to_signed(-5, 8),
    to_signed(-5, 8),
    to_signed(-6, 8),
    to_signed(-7, 8),
    to_signed(-6, 8),
    to_signed(-4, 8),
    to_signed(-1, 8),
    to_signed(-1, 8),
    to_signed(-2, 8),
    to_signed(-3, 8),
    to_signed(-2, 8),
    to_signed(-2, 8),
    to_signed(-2, 8),
    to_signed(-2, 8),
    to_signed(0, 8),
    to_signed(1, 8),
    to_signed(1, 8),
    to_signed(1, 8),
    to_signed(1, 8),
    to_signed(1, 8),
    to_signed(2, 8),
    to_signed(3, 8),
    to_signed(4, 8),
    to_signed(5, 8),
    to_signed(7, 8),
    to_signed(8, 8),
    to_signed(9, 8),
    to_signed(11, 8),
    to_signed(12, 8),
    to_signed(13, 8),
    to_signed(14, 8),
    to_signed(14, 8),
    to_signed(13, 8),
    to_signed(11, 8),
    to_signed(10, 8),
    to_signed(10, 8),
    to_signed(9, 8),
    to_signed(9, 8),
    to_signed(7, 8),
    to_signed(5, 8),
    to_signed(4, 8),
    to_signed(3, 8),
    to_signed(3, 8),
    to_signed(2, 8),
    to_signed(2, 8),
    to_signed(1, 8),
    to_signed(0, 8),
    to_signed(-2, 8),
    to_signed(-3, 8),
    to_signed(-2, 8),
    to_signed(-1, 8),
    to_signed(-1, 8),
    to_signed(-1, 8),
    to_signed(-2, 8),
    to_signed(-4, 8),
    to_signed(-7, 8),
    to_signed(-9, 8),
    to_signed(-11, 8),
    to_signed(-12, 8),
    to_signed(-12, 8),
    to_signed(-12, 8),
    to_signed(-12, 8),
    to_signed(-13, 8),
    to_signed(-12, 8),
    to_signed(-12, 8),
    to_signed(-11, 8),
    to_signed(-11, 8),
    to_signed(-11, 8),
    to_signed(-11, 8),
    to_signed(-9, 8),
    to_signed(-8, 8),
    to_signed(-7, 8),
    to_signed(-7, 8),
    to_signed(-6, 8),
    to_signed(-5, 8),
    to_signed(-5, 8),
    to_signed(-5, 8),
    to_signed(-6, 8),
    to_signed(-5, 8),
    to_signed(-4, 8),
    to_signed(-4, 8),
    to_signed(-4, 8),
    to_signed(-5, 8),
    to_signed(-5, 8),
    to_signed(-4, 8),
    to_signed(-3, 8),
    to_signed(-2, 8),
    to_signed(-1, 8),
    to_signed(-1, 8),
    to_signed(-1, 8),
    to_signed(-1, 8),
    to_signed(-1, 8),
    to_signed(1, 8),
    to_signed(3, 8),
    to_signed(6, 8),
    to_signed(8, 8),
    to_signed(9, 8),
    to_signed(8, 8),
    to_signed(8, 8),
    to_signed(8, 8),
    to_signed(8, 8),
    to_signed(8, 8),
    to_signed(8, 8),
    to_signed(9, 8),
    to_signed(8, 8),
    to_signed(7, 8),
    to_signed(4, 8),
    to_signed(3, 8),
    to_signed(2, 8),
    to_signed(3, 8),
    to_signed(3, 8),
    to_signed(4, 8),
    to_signed(3, 8),
    to_signed(2, 8),
    to_signed(0, 8),
    to_signed(0, 8),
    to_signed(0, 8),
    to_signed(1, 8),
    to_signed(1, 8),
    to_signed(1, 8),
    to_signed(-1, 8),
    to_signed(-3, 8),
    to_signed(-4, 8),
    to_signed(-5, 8),
    to_signed(-6, 8),
    to_signed(-7, 8),
    to_signed(-9, 8),
    to_signed(-9, 8),
    to_signed(-8, 8),
    to_signed(-7, 8),
    to_signed(-6, 8),
    to_signed(-6, 8),
    to_signed(-6, 8),
    to_signed(-6, 8),
    to_signed(-6, 8),
    to_signed(-5, 8),
    to_signed(-5, 8),
    to_signed(-4, 8),
    to_signed(-2, 8),
    to_signed(-1, 8),
    to_signed(1, 8),
    to_signed(2, 8),
    to_signed(2, 8),
    to_signed(1, 8),
    to_signed(0, 8),
    to_signed(-1, 8),
    to_signed(-2, 8),
    to_signed(-3, 8),
    to_signed(-3, 8),
    to_signed(-2, 8),
    to_signed(-2, 8),
    to_signed(-1, 8),
    to_signed(-1, 8),
    to_signed(0, 8),
    to_signed(0, 8),
    to_signed(1, 8),
    to_signed(0, 8),
    to_signed(0, 8),
    to_signed(1, 8),
    to_signed(3, 8),
    to_signed(5, 8),
    to_signed(7, 8),
    to_signed(7, 8),
    to_signed(6, 8),
    to_signed(4, 8),
    to_signed(3, 8),
    to_signed(2, 8),
    to_signed(1, 8),
    to_signed(0, 8),
    to_signed(0, 8),
    to_signed(0, 8),
    to_signed(0, 8),
    to_signed(-1, 8),
    to_signed(-2, 8),
    to_signed(-3, 8),
    to_signed(-2, 8),
    to_signed(-2, 8),
    to_signed(-2, 8),
    to_signed(-2, 8),
    to_signed(-3, 8),
    to_signed(-3, 8),
    to_signed(-4, 8),
    to_signed(-3, 8),
    to_signed(-2, 8),
    to_signed(-1, 8),
    to_signed(0, 8),
    to_signed(-1, 8),
    to_signed(-3, 8),
    to_signed(-5, 8),
    to_signed(-6, 8),
    to_signed(-5, 8),
    to_signed(-4, 8),
    to_signed(-3, 8),
    to_signed(-1, 8),
    to_signed(0, 8),
    to_signed(0, 8),
    to_signed(0, 8),
    to_signed(-1, 8),
    to_signed(0, 8),
    to_signed(0, 8),
    to_signed(1, 8),
    to_signed(1, 8),
    to_signed(2, 8),
    to_signed(3, 8),
    to_signed(4, 8),
    to_signed(6, 8),
    to_signed(7, 8),
    to_signed(8, 8),
    to_signed(8, 8),
    to_signed(8, 8),
    to_signed(7, 8),
    to_signed(6, 8),
    to_signed(6, 8),
    to_signed(5, 8),
    to_signed(4, 8),
    to_signed(3, 8),
    to_signed(2, 8),
    to_signed(1, 8),
    to_signed(1, 8),
    to_signed(1, 8),
    to_signed(1, 8),
    to_signed(1, 8),
    to_signed(0, 8),
    to_signed(0, 8),
    to_signed(-1, 8),
    to_signed(-1, 8),
    to_signed(0, 8),
    to_signed(1, 8),
    to_signed(1, 8),
    to_signed(0, 8),
    to_signed(-1, 8),
    to_signed(-2, 8),
    to_signed(-5, 8),
    to_signed(-6, 8),
    to_signed(-7, 8),
    to_signed(-8, 8),
    to_signed(-9, 8),
    to_signed(-10, 8),
    to_signed(-10, 8),
    to_signed(-10, 8),
    to_signed(-9, 8),
    to_signed(-9, 8),
    to_signed(-10, 8),
    to_signed(-10, 8),
    to_signed(-10, 8),
    to_signed(-10, 8),
    to_signed(-10, 8),
    to_signed(-9, 8),
    to_signed(-8, 8),
    to_signed(-7, 8),
    to_signed(-7, 8),
    to_signed(-8, 8),
    to_signed(-8, 8),
    to_signed(-8, 8),
    to_signed(-7, 8),
    to_signed(-7, 8),
    to_signed(-8, 8),
    to_signed(-8, 8),
    to_signed(-8, 8),
    to_signed(-8, 8),
    to_signed(-7, 8),
    to_signed(-6, 8),
    to_signed(-5, 8),
    to_signed(-4, 8),
    to_signed(-2, 8),
    to_signed(-1, 8),
    to_signed(0, 8),
    to_signed(1, 8),
    to_signed(2, 8),
    to_signed(3, 8),
    to_signed(4, 8),
    to_signed(5, 8),
    to_signed(8, 8),
    to_signed(9, 8),
    to_signed(10, 8),
    to_signed(9, 8),
    to_signed(7, 8),
    to_signed(6, 8),
    to_signed(5, 8),
    to_signed(4, 8),
    to_signed(3, 8),
    to_signed(2, 8),
    to_signed(2, 8),
    to_signed(1, 8),
    to_signed(1, 8),
    to_signed(0, 8),
    to_signed(-1, 8),
    to_signed(-1, 8),
    to_signed(-1, 8),
    to_signed(-1, 8),
    to_signed(-2, 8),
    to_signed(-2, 8),
    to_signed(-2, 8),
    to_signed(-2, 8),
    to_signed(-1, 8),
    to_signed(-1, 8),
    to_signed(-2, 8),
    to_signed(-4, 8),
    to_signed(-6, 8),
    to_signed(-8, 8),
    to_signed(-10, 8),
    to_signed(-11, 8),
    to_signed(-12, 8),
    to_signed(-12, 8),
    to_signed(-11, 8),
    to_signed(-11, 8),
    to_signed(-11, 8),
    to_signed(-10, 8),
    to_signed(-10, 8),
    to_signed(-9, 8),
    to_signed(-9, 8),
    to_signed(-8, 8),
    to_signed(-8, 8),
    to_signed(-7, 8),
    to_signed(-6, 8),
    to_signed(-3, 8),
    to_signed(-2, 8),
    to_signed(-1, 8),
    to_signed(-2, 8),
    to_signed(-2, 8),
    to_signed(-2, 8),
    to_signed(-1, 8),
    to_signed(0, 8),
    to_signed(1, 8),
    to_signed(2, 8),
    to_signed(2, 8),
    to_signed(3, 8),
    to_signed(4, 8),
    to_signed(5, 8),
    to_signed(6, 8),
    to_signed(8, 8),
    to_signed(9, 8),
    to_signed(11, 8),
    to_signed(12, 8),
    to_signed(12, 8),
    to_signed(13, 8),
    to_signed(13, 8),
    to_signed(14, 8),
    to_signed(15, 8),
    to_signed(15, 8),
    to_signed(14, 8),
    to_signed(13, 8),
    to_signed(12, 8),
    to_signed(11, 8),
    to_signed(9, 8),
    to_signed(7, 8),
    to_signed(5, 8),
    to_signed(4, 8),
    to_signed(3, 8),
    to_signed(2, 8),
    to_signed(2, 8),
    to_signed(1, 8),
    to_signed(0, 8),
    to_signed(-1, 8),
    to_signed(-2, 8),
    to_signed(-3, 8),
    to_signed(-4, 8),
    to_signed(-4, 8),
    to_signed(-3, 8),
    to_signed(-2, 8),
    to_signed(-1, 8),
    to_signed(-2, 8),
    to_signed(-3, 8),
    to_signed(-5, 8),
    to_signed(-6, 8),
    to_signed(-6, 8),
    to_signed(-7, 8),
    to_signed(-8, 8),
    to_signed(-8, 8),
    to_signed(-9, 8),
    to_signed(-9, 8),
    to_signed(-8, 8),
    to_signed(-6, 8),
    to_signed(-5, 8),
    to_signed(-3, 8),
    to_signed(-2, 8),
    to_signed(0, 8),
    to_signed(0, 8),
    to_signed(1, 8),
    to_signed(2, 8),
    to_signed(2, 8),
    to_signed(4, 8),
    to_signed(5, 8),
    to_signed(5, 8),
    to_signed(5, 8),
    to_signed(4, 8),
    to_signed(5, 8),
    to_signed(6, 8),
    to_signed(6, 8),
    to_signed(6, 8),
    to_signed(6, 8),
    to_signed(7, 8),
    to_signed(8, 8),
    to_signed(9, 8),
    to_signed(10, 8),
    to_signed(10, 8),
    to_signed(10, 8),
    to_signed(9, 8),
    to_signed(9, 8),
    to_signed(8, 8),
    to_signed(8, 8),
    to_signed(8, 8),
    to_signed(9, 8),
    to_signed(10, 8),
    to_signed(10, 8),
    to_signed(9, 8),
    to_signed(8, 8),
    to_signed(8, 8),
    to_signed(7, 8),
    to_signed(6, 8),
    to_signed(5, 8),
    to_signed(4, 8),
    to_signed(3, 8),
    to_signed(2, 8),
    to_signed(0, 8),
    to_signed(-2, 8),
    to_signed(-3, 8),
    to_signed(-4, 8),
    to_signed(-4, 8),
    to_signed(-5, 8),
    to_signed(-6, 8),
    to_signed(-5, 8),
    to_signed(-5, 8),
    to_signed(-5, 8),
    to_signed(-6, 8),
    to_signed(-5, 8),
    to_signed(-5, 8),
    to_signed(-5, 8),
    to_signed(-7, 8),
    to_signed(-8, 8),
    to_signed(-8, 8),
    to_signed(-8, 8),
    to_signed(-8, 8),
    to_signed(-9, 8),
    to_signed(-10, 8),
    to_signed(-10, 8),
    to_signed(-9, 8),
    to_signed(-10, 8),
    to_signed(-9, 8),
    to_signed(-8, 8),
    to_signed(-7, 8),
    to_signed(-6, 8),
    to_signed(-5, 8),
    to_signed(-4, 8),
    to_signed(-2, 8),
    to_signed(-1, 8),
    to_signed(-1, 8),
    to_signed(0, 8),
    to_signed(1, 8),
    to_signed(3, 8),
    to_signed(4, 8),
    to_signed(4, 8),
    to_signed(4, 8),
    to_signed(4, 8),
    to_signed(3, 8),
    to_signed(3, 8),
    to_signed(3, 8),
    to_signed(2, 8),
    to_signed(3, 8),
    to_signed(4, 8),
    to_signed(4, 8),
    to_signed(4, 8),
    to_signed(4, 8),
    to_signed(4, 8),
    to_signed(5, 8),
    to_signed(5, 8),
    to_signed(6, 8),
    to_signed(8, 8),
    to_signed(9, 8),
    to_signed(8, 8),
    to_signed(7, 8),
    to_signed(6, 8),
    to_signed(5, 8),
    to_signed(3, 8),
    to_signed(2, 8),
    to_signed(1, 8),
    to_signed(0, 8),
    to_signed(0, 8),
    to_signed(-1, 8),
    to_signed(-2, 8),
    to_signed(-3, 8),
    to_signed(-4, 8),
    to_signed(-4, 8),
    to_signed(-3, 8),
    to_signed(-3, 8),
    to_signed(-2, 8),
    to_signed(-3, 8),
    to_signed(-4, 8),
    to_signed(-6, 8),
    to_signed(-7, 8),
    to_signed(-7, 8),
    to_signed(-6, 8),
    to_signed(-5, 8),
    to_signed(-4, 8),
    to_signed(-5, 8),
    to_signed(-6, 8),
    to_signed(-7, 8),
    to_signed(-8, 8),
    to_signed(-9, 8),
    to_signed(-8, 8),
    to_signed(-6, 8),
    to_signed(-6, 8),
    to_signed(-6, 8),
    to_signed(-6, 8),
    to_signed(-6, 8),
    to_signed(-5, 8),
    to_signed(-4, 8),
    to_signed(-2, 8),
    to_signed(-1, 8),
    to_signed(1, 8),
    to_signed(1, 8),
    to_signed(1, 8),
    to_signed(1, 8),
    to_signed(2, 8),
    to_signed(2, 8),
    to_signed(3, 8),
    to_signed(4, 8),
    to_signed(4, 8),
    to_signed(4, 8),
    to_signed(3, 8),
    to_signed(3, 8),
    to_signed(2, 8),
    to_signed(1, 8),
    to_signed(0, 8),
    to_signed(0, 8),
    to_signed(1, 8),
    to_signed(1, 8),
    to_signed(2, 8),
    to_signed(3, 8),
    to_signed(3, 8),
    to_signed(3, 8),
    to_signed(3, 8),
    to_signed(2, 8),
    to_signed(1, 8),
    to_signed(0, 8),
    to_signed(1, 8),
    to_signed(2, 8),
    to_signed(3, 8),
    to_signed(3, 8),
    to_signed(2, 8),
    to_signed(2, 8),
    to_signed(1, 8),
    to_signed(0, 8),
    to_signed(0, 8),
    to_signed(-1, 8),
    to_signed(-1, 8),
    to_signed(-2, 8),
    to_signed(-3, 8),
    to_signed(-4, 8),
    to_signed(-3, 8),
    to_signed(-2, 8),
    to_signed(-1, 8),
    to_signed(-1, 8),
    to_signed(-1, 8),
    to_signed(-1, 8),
    to_signed(-2, 8),
    to_signed(-2, 8),
    to_signed(-2, 8),
    to_signed(-2, 8),
    to_signed(-2, 8),
    to_signed(-2, 8),
    to_signed(-2, 8),
    to_signed(-1, 8),
    to_signed(-1, 8),
    to_signed(-3, 8),
    to_signed(-4, 8),
    to_signed(-5, 8),
    to_signed(-6, 8),
    to_signed(-7, 8),
    to_signed(-8, 8),
    to_signed(-8, 8),
    to_signed(-7, 8),
    to_signed(-5, 8),
    to_signed(-5, 8),
    to_signed(-4, 8),
    to_signed(-5, 8),
    to_signed(-5, 8),
    to_signed(-6, 8),
    to_signed(-5, 8),
    to_signed(-4, 8),
    to_signed(-3, 8),
    to_signed(-2, 8),
    to_signed(-2, 8),
    to_signed(-3, 8),
    to_signed(-5, 8),
    to_signed(-6, 8),
    to_signed(-6, 8),
    to_signed(-6, 8),
    to_signed(-5, 8),
    to_signed(-5, 8),
    to_signed(-5, 8),
    to_signed(-5, 8),
    to_signed(-5, 8),
    to_signed(-5, 8),
    to_signed(-5, 8),
    to_signed(-4, 8),
    to_signed(-4, 8),
    to_signed(-4, 8),
    to_signed(-6, 8),
    to_signed(-6, 8),
    to_signed(-4, 8),
    to_signed(-2, 8),
    to_signed(-2, 8),
    to_signed(-1, 8),
    to_signed(-1, 8),
    to_signed(-1, 8),
    to_signed(-2, 8),
    to_signed(-3, 8),
    to_signed(-3, 8),
    to_signed(-3, 8),
    to_signed(-3, 8),
    to_signed(-3, 8),
    to_signed(-3, 8),
    to_signed(-3, 8),
    to_signed(-3, 8),
    to_signed(-3, 8),
    to_signed(-1, 8),
    to_signed(0, 8),
    to_signed(0, 8),
    to_signed(0, 8),
    to_signed(-1, 8),
    to_signed(-1, 8),
    to_signed(0, 8),
    to_signed(2, 8),
    to_signed(3, 8),
    to_signed(4, 8),
    to_signed(4, 8),
    to_signed(3, 8),
    to_signed(1, 8),
    to_signed(-1, 8),
    to_signed(-2, 8),
    to_signed(-2, 8),
    to_signed(-2, 8),
    to_signed(-2, 8),
    to_signed(-2, 8),
    to_signed(-1, 8),
    to_signed(-1, 8),
    to_signed(-1, 8),
    to_signed(0, 8),
    to_signed(1, 8),
    to_signed(1, 8),
    to_signed(0, 8),
    to_signed(0, 8),
    to_signed(0, 8),
    to_signed(1, 8),
    to_signed(1, 8),
    to_signed(1, 8),
    to_signed(1, 8),
    to_signed(1, 8),
    to_signed(1, 8),
    to_signed(-1, 8),
    to_signed(-1, 8),
    to_signed(-2, 8),
    to_signed(-3, 8),
    to_signed(-4, 8),
    to_signed(-5, 8),
    to_signed(-5, 8),
    to_signed(-5, 8),
    to_signed(-5, 8),
    to_signed(-5, 8),
    to_signed(-5, 8),
    to_signed(-4, 8),
    to_signed(-4, 8),
    to_signed(-4, 8),
    to_signed(-4, 8),
    to_signed(-3, 8),
    to_signed(-2, 8),
    to_signed(-2, 8),
    to_signed(-1, 8),
    to_signed(-1, 8),
    to_signed(0, 8),
    to_signed(-1, 8),
    to_signed(-1, 8),
    to_signed(-1, 8),
    to_signed(0, 8),
    to_signed(-1, 8),
    to_signed(-3, 8),
    to_signed(-4, 8),
    to_signed(-4, 8),
    to_signed(-2, 8),
    to_signed(0, 8),
    to_signed(2, 8),
    to_signed(4, 8),
    to_signed(5, 8),
    to_signed(5, 8),
    to_signed(5, 8),
    to_signed(5, 8),
    to_signed(6, 8),
    to_signed(8, 8),
    to_signed(10, 8),
    to_signed(10, 8),
    to_signed(10, 8),
    to_signed(9, 8),
    to_signed(9, 8),
    to_signed(9, 8),
    to_signed(7, 8),
    to_signed(6, 8),
    to_signed(4, 8),
    to_signed(3, 8),
    to_signed(3, 8),
    to_signed(3, 8),
    to_signed(3, 8),
    to_signed(4, 8),
    to_signed(5, 8),
    to_signed(5, 8),
    to_signed(3, 8),
    to_signed(2, 8),
    to_signed(1, 8),
    to_signed(1, 8),
    to_signed(1, 8),
    to_signed(1, 8),
    to_signed(2, 8),
    to_signed(2, 8),
    to_signed(2, 8),
    to_signed(1, 8),
    to_signed(0, 8),
    to_signed(-1, 8),
    to_signed(-2, 8),
    to_signed(-3, 8),
    to_signed(-5, 8),
    to_signed(-7, 8),
    to_signed(-7, 8),
    to_signed(-7, 8),
    to_signed(-6, 8),
    to_signed(-6, 8),
    to_signed(-5, 8),
    to_signed(-4, 8),
    to_signed(-4, 8),
    to_signed(-5, 8),
    to_signed(-5, 8),
    to_signed(-4, 8),
    to_signed(-3, 8),
    to_signed(-2, 8),
    to_signed(-2, 8),
    to_signed(-1, 8),
    to_signed(1, 8),
    to_signed(1, 8),
    to_signed(1, 8),
    to_signed(1, 8),
    to_signed(1, 8),
    to_signed(-1, 8),
    to_signed(-2, 8),
    to_signed(-2, 8),
    to_signed(-1, 8),
    to_signed(1, 8),
    to_signed(3, 8),
    to_signed(4, 8),
    to_signed(5, 8),
    to_signed(5, 8),
    to_signed(4, 8),
    to_signed(4, 8),
    to_signed(6, 8),
    to_signed(8, 8),
    to_signed(8, 8),
    to_signed(8, 8),
    to_signed(8, 8),
    to_signed(8, 8),
    to_signed(8, 8),
    to_signed(8, 8),
    to_signed(7, 8),
    to_signed(6, 8),
    to_signed(5, 8),
    to_signed(4, 8),
    to_signed(3, 8),
    to_signed(3, 8),
    to_signed(2, 8),
    to_signed(1, 8),
    to_signed(0, 8),
    to_signed(0, 8),
    to_signed(0, 8),
    to_signed(1, 8),
    to_signed(1, 8),
    to_signed(1, 8),
    to_signed(1, 8),
    to_signed(1, 8),
    to_signed(1, 8),
    to_signed(0, 8),
    to_signed(0, 8),
    to_signed(0, 8),
    to_signed(1, 8),
    to_signed(1, 8),
    to_signed(1, 8),
    to_signed(1, 8),
    to_signed(1, 8),
    to_signed(1, 8),
    to_signed(0, 8),
    to_signed(0, 8),
    to_signed(-1, 8),
    to_signed(-1, 8),
    to_signed(-2, 8),
    to_signed(-1, 8),
    to_signed(0, 8),
    to_signed(1, 8),
    to_signed(2, 8),
    to_signed(4, 8),
    to_signed(4, 8),
    to_signed(4, 8),
    to_signed(4, 8),
    to_signed(6, 8),
    to_signed(8, 8),
    to_signed(10, 8),
    to_signed(10, 8),
    to_signed(10, 8),
    to_signed(9, 8),
    to_signed(7, 8),
    to_signed(5, 8),
    to_signed(5, 8),
    to_signed(5, 8),
    to_signed(4, 8),
    to_signed(3, 8),
    to_signed(2, 8),
    to_signed(3, 8),
    to_signed(4, 8),
    to_signed(5, 8),
    to_signed(5, 8),
    to_signed(7, 8),
    to_signed(8, 8),
    to_signed(7, 8),
    to_signed(6, 8),
    to_signed(6, 8),
    to_signed(6, 8),
    to_signed(6, 8),
    to_signed(5, 8),
    to_signed(4, 8),
    to_signed(4, 8),
    to_signed(3, 8),
    to_signed(2, 8),
    to_signed(0, 8),
    to_signed(-1, 8),
    to_signed(-2, 8),
    to_signed(-3, 8),
    to_signed(-5, 8),
    to_signed(-5, 8),
    to_signed(-6, 8),
    to_signed(-6, 8),
    to_signed(-6, 8),
    to_signed(-5, 8),
    to_signed(-4, 8),
    to_signed(-4, 8),
    to_signed(-5, 8),
    to_signed(-6, 8),
    to_signed(-6, 8),
    to_signed(-7, 8),
    to_signed(-7, 8),
    to_signed(-6, 8),
    to_signed(-5, 8),
    to_signed(-4, 8),
    to_signed(-4, 8),
    to_signed(-4, 8),
    to_signed(-4, 8),
    to_signed(-5, 8),
    to_signed(-6, 8),
    to_signed(-7, 8),
    to_signed(-6, 8),
    to_signed(-5, 8),
    to_signed(-4, 8),
    to_signed(-3, 8),
    to_signed(-2, 8),
    to_signed(1, 8),
    to_signed(2, 8),
    to_signed(2, 8),
    to_signed(2, 8),
    to_signed(2, 8),
    to_signed(3, 8),
    to_signed(3, 8),
    to_signed(3, 8),
    to_signed(3, 8),
    to_signed(4, 8),
    to_signed(5, 8),
    to_signed(6, 8),
    to_signed(5, 8),
    to_signed(4, 8),
    to_signed(3, 8),
    to_signed(1, 8),
    to_signed(-1, 8),
    to_signed(-2, 8),
    to_signed(-2, 8),
    to_signed(-1, 8),
    to_signed(-1, 8),
    to_signed(-1, 8),
    to_signed(-1, 8),
    to_signed(-1, 8),
    to_signed(-1, 8),
    to_signed(-1, 8),
    to_signed(-1, 8),
    to_signed(-1, 8),
    to_signed(-1, 8),
    to_signed(-2, 8),
    to_signed(-2, 8),
    to_signed(-2, 8),
    to_signed(-3, 8),
    to_signed(-4, 8),
    to_signed(-4, 8),
    to_signed(-5, 8),
    to_signed(-6, 8),
    to_signed(-7, 8),
    to_signed(-8, 8),
    to_signed(-9, 8),
    to_signed(-8, 8),
    to_signed(-7, 8),
    to_signed(-6, 8),
    to_signed(-4, 8),
    to_signed(-2, 8),
    to_signed(-1, 8),
    to_signed(-2, 8),
    to_signed(-4, 8),
    to_signed(-5, 8),
    to_signed(-5, 8),
    to_signed(-3, 8),
    to_signed(-1, 8),
    to_signed(1, 8),
    to_signed(2, 8),
    to_signed(2, 8),
    to_signed(2, 8),
    to_signed(1, 8),
    to_signed(1, 8),
    to_signed(1, 8),
    to_signed(0, 8),
    to_signed(-2, 8),
    to_signed(-2, 8),
    to_signed(-1, 8),
    to_signed(1, 8),
    to_signed(2, 8),
    to_signed(3, 8),
    to_signed(3, 8),
    to_signed(2, 8),
    to_signed(2, 8),
    to_signed(2, 8),
    to_signed(3, 8),
    to_signed(5, 8),
    to_signed(6, 8),
    to_signed(6, 8),
    to_signed(5, 8),
    to_signed(4, 8),
    to_signed(2, 8),
    to_signed(0, 8),
    to_signed(-1, 8),
    to_signed(-1, 8),
    to_signed(-1, 8),
    to_signed(-2, 8),
    to_signed(-3, 8),
    to_signed(-4, 8),
    to_signed(-4, 8),
    to_signed(-5, 8),
    to_signed(-6, 8),
    to_signed(-6, 8),
    to_signed(-6, 8),
    to_signed(-5, 8),
    to_signed(-4, 8),
    to_signed(-3, 8),
    to_signed(-2, 8),
    to_signed(-2, 8),
    to_signed(-3, 8),
    to_signed(-4, 8),
    to_signed(-5, 8),
    to_signed(-5, 8),
    to_signed(-6, 8),
    to_signed(-6, 8),
    to_signed(-4, 8),
    to_signed(-4, 8),
    to_signed(-5, 8),
    to_signed(-8, 8),
    to_signed(-9, 8),
    to_signed(-8, 8),
    to_signed(-6, 8),
    to_signed(-4, 8),
    to_signed(-4, 8),
    to_signed(-3, 8),
    to_signed(-4, 8),
    to_signed(-4, 8),
    to_signed(-3, 8),
    to_signed(-2, 8),
    to_signed(-1, 8),
    to_signed(0, 8),
    to_signed(1, 8),
    to_signed(3, 8),
    to_signed(3, 8),
    to_signed(2, 8),
    to_signed(1, 8),
    to_signed(1, 8),
    to_signed(0, 8),
    to_signed(-2, 8),
    to_signed(-3, 8),
    to_signed(-3, 8),
    to_signed(-2, 8),
    to_signed(-1, 8),
    to_signed(-1, 8),
    to_signed(-1, 8),
    to_signed(-1, 8),
    to_signed(-1, 8),
    to_signed(-1, 8),
    to_signed(0, 8),
    to_signed(1, 8),
    to_signed(3, 8),
    to_signed(4, 8),
    to_signed(4, 8),
    to_signed(3, 8),
    to_signed(1, 8),
    to_signed(0, 8),
    to_signed(0, 8),
    to_signed(1, 8),
    to_signed(1, 8),
    to_signed(0, 8),
    to_signed(-1, 8),
    to_signed(-2, 8),
    to_signed(-4, 8),
    to_signed(-5, 8),
    to_signed(-6, 8),
    to_signed(-7, 8),
    to_signed(-6, 8),
    to_signed(-5, 8),
    to_signed(-4, 8),
    to_signed(-4, 8),
    to_signed(-3, 8),
    to_signed(-3, 8),
    to_signed(-3, 8),
    to_signed(-4, 8),
    to_signed(-4, 8),
    to_signed(-4, 8),
    to_signed(-3, 8),
    to_signed(-3, 8),
    to_signed(-3, 8),
    to_signed(-3, 8),
    to_signed(-2, 8),
    to_signed(-2, 8),
    to_signed(-3, 8),
    to_signed(-5, 8),
    to_signed(-7, 8),
    to_signed(-8, 8),
    to_signed(-8, 8),
    to_signed(-7, 8),
    to_signed(-4, 8),
    to_signed(-2, 8),
    to_signed(-1, 8),
    to_signed(-1, 8),
    to_signed(-1, 8),
    to_signed(-1, 8),
    to_signed(-1, 8),
    to_signed(-1, 8),
    to_signed(-1, 8),
    to_signed(0, 8),
    to_signed(1, 8),
    to_signed(1, 8),
    to_signed(2, 8),
    to_signed(2, 8),
    to_signed(1, 8),
    to_signed(-1, 8),
    to_signed(-2, 8),
    to_signed(-2, 8),
    to_signed(-2, 8),
    to_signed(-3, 8),
    to_signed(-3, 8),
    to_signed(-2, 8),
    to_signed(-1, 8),
    to_signed(0, 8),
    to_signed(1, 8),
    to_signed(2, 8),
    to_signed(1, 8),
    to_signed(0, 8),
    to_signed(0, 8),
    to_signed(1, 8),
    to_signed(1, 8),
    to_signed(1, 8),
    to_signed(0, 8),
    to_signed(1, 8),
    to_signed(1, 8),
    to_signed(0, 8),
    to_signed(-1, 8),
    to_signed(-2, 8),
    to_signed(-2, 8),
    to_signed(-4, 8),
    to_signed(-6, 8),
    to_signed(-7, 8),
    to_signed(-7, 8),
    to_signed(-6, 8),
    to_signed(-4, 8),
    to_signed(-3, 8),
    to_signed(-1, 8),
    to_signed(-1, 8),
    to_signed(-2, 8),
    to_signed(-2, 8),
    to_signed(-2, 8),
    to_signed(-2, 8),
    to_signed(-3, 8),
    to_signed(-3, 8),
    to_signed(-2, 8),
    to_signed(-1, 8),
    to_signed(-1, 8),
    to_signed(-2, 8),
    to_signed(-3, 8),
    to_signed(-4, 8),
    to_signed(-4, 8),
    to_signed(-4, 8),
    to_signed(-4, 8),
    to_signed(-3, 8),
    to_signed(-2, 8),
    to_signed(0, 8),
    to_signed(1, 8),
    to_signed(0, 8),
    to_signed(-2, 8),
    to_signed(-2, 8),
    to_signed(-2, 8),
    to_signed(0, 8),
    to_signed(1, 8),
    to_signed(2, 8),
    to_signed(3, 8),
    to_signed(4, 8),
    to_signed(4, 8),
    to_signed(2, 8),
    to_signed(2, 8),
    to_signed(2, 8),
    to_signed(2, 8),
    to_signed(2, 8),
    to_signed(3, 8),
    to_signed(3, 8),
    to_signed(3, 8),
    to_signed(4, 8),
    to_signed(4, 8),
    to_signed(4, 8),
    to_signed(4, 8),
    to_signed(4, 8),
    to_signed(4, 8),
    to_signed(4, 8),
    to_signed(4, 8),
    to_signed(3, 8),
    to_signed(3, 8),
    to_signed(3, 8),
    to_signed(3, 8),
    to_signed(4, 8),
    to_signed(4, 8),
    to_signed(4, 8),
    to_signed(3, 8),
    to_signed(3, 8),
    to_signed(2, 8),
    to_signed(1, 8),
    to_signed(-1, 8),
    to_signed(-2, 8),
    to_signed(-3, 8),
    to_signed(-2, 8),
    to_signed(-1, 8),
    to_signed(-1, 8),
    to_signed(0, 8),
    to_signed(-1, 8),
    to_signed(-3, 8),
    to_signed(-4, 8),
    to_signed(-5, 8),
    to_signed(-5, 8),
    to_signed(-4, 8),
    to_signed(-2, 8),
    to_signed(-1, 8),
    to_signed(-1, 8),
    to_signed(-2, 8),
    to_signed(-3, 8),
    to_signed(-4, 8),
    to_signed(-4, 8),
    to_signed(-6, 8),
    to_signed(-6, 8),
    to_signed(-6, 8),
    to_signed(-4, 8),
    to_signed(-5, 8),
    to_signed(-6, 8),
    to_signed(-7, 8),
    to_signed(-7, 8),
    to_signed(-6, 8),
    to_signed(-5, 8),
    to_signed(-5, 8),
    to_signed(-4, 8),
    to_signed(-4, 8),
    to_signed(-4, 8),
    to_signed(-3, 8),
    to_signed(-1, 8),
    to_signed(-2, 8),
    to_signed(-3, 8),
    to_signed(-3, 8),
    to_signed(-2, 8),
    to_signed(-1, 8),
    to_signed(0, 8),
    to_signed(1, 8),
    to_signed(3, 8),
    to_signed(3, 8),
    to_signed(0, 8),
    to_signed(-3, 8),
    to_signed(-3, 8),
    to_signed(-1, 8),
    to_signed(0, 8),
    to_signed(2, 8),
    to_signed(3, 8),
    to_signed(5, 8),
    to_signed(5, 8),
    to_signed(3, 8),
    to_signed(1, 8),
    to_signed(0, 8),
    to_signed(-1, 8),
    to_signed(-1, 8),
    to_signed(1, 8),
    to_signed(3, 8),
    to_signed(5, 8),
    to_signed(5, 8),
    to_signed(5, 8),
    to_signed(3, 8),
    to_signed(0, 8),
    to_signed(-3, 8),
    to_signed(-5, 8),
    to_signed(-6, 8),
    to_signed(-6, 8),
    to_signed(-6, 8),
    to_signed(-5, 8),
    to_signed(-3, 8),
    to_signed(-1, 8),
    to_signed(-2, 8),
    to_signed(-3, 8),
    to_signed(-5, 8),
    to_signed(-6, 8),
    to_signed(-6, 8),
    to_signed(-6, 8),
    to_signed(-7, 8),
    to_signed(-6, 8),
    to_signed(-6, 8),
    to_signed(-5, 8),
    to_signed(-6, 8),
    to_signed(-6, 8),
    to_signed(-6, 8),
    to_signed(-5, 8),
    to_signed(-6, 8),
    to_signed(-8, 8),
    to_signed(-10, 8),
    to_signed(-10, 8),
    to_signed(-9, 8),
    to_signed(-8, 8),
    to_signed(-7, 8),
    to_signed(-5, 8),
    to_signed(-3, 8),
    to_signed(-2, 8),
    to_signed(-2, 8),
    to_signed(-4, 8),
    to_signed(-5, 8),
    to_signed(-5, 8),
    to_signed(-6, 8),
    to_signed(-5, 8),
    to_signed(-2, 8),
    to_signed(0, 8),
    to_signed(2, 8),
    to_signed(2, 8),
    to_signed(0, 8),
    to_signed(-2, 8),
    to_signed(-3, 8),
    to_signed(-3, 8),
    to_signed(-3, 8),
    to_signed(-4, 8),
    to_signed(-3, 8),
    to_signed(-2, 8),
    to_signed(-1, 8),
    to_signed(-1, 8),
    to_signed(-1, 8),
    to_signed(-1, 8),
    to_signed(-1, 8),
    to_signed(-1, 8),
    to_signed(-1, 8),
    to_signed(-1, 8),
    to_signed(0, 8),
    to_signed(2, 8),
    to_signed(2, 8),
    to_signed(2, 8),
    to_signed(1, 8),
    to_signed(1, 8),
    to_signed(1, 8),
    to_signed(1, 8),
    to_signed(2, 8),
    to_signed(1, 8),
    to_signed(0, 8),
    to_signed(0, 8),
    to_signed(0, 8),
    to_signed(-1, 8),
    to_signed(-2, 8),
    to_signed(-2, 8),
    to_signed(1, 8),
    to_signed(3, 8),
    to_signed(2, 8),
    to_signed(1, 8),
    to_signed(1, 8),
    to_signed(2, 8),
    to_signed(2, 8),
    to_signed(0, 8),
    to_signed(-1, 8),
    to_signed(0, 8),
    to_signed(2, 8),
    to_signed(2, 8),
    to_signed(1, 8),
    to_signed(0, 8),
    to_signed(-1, 8),
    to_signed(-2, 8),
    to_signed(-3, 8),
    to_signed(-3, 8),
    to_signed(-3, 8),
    to_signed(-3, 8),
    to_signed(-2, 8),
    to_signed(-2, 8),
    to_signed(-3, 8),
    to_signed(-3, 8),
    to_signed(-2, 8),
    to_signed(-1, 8),
    to_signed(1, 8),
    to_signed(1, 8),
    to_signed(2, 8),
    to_signed(2, 8),
    to_signed(3, 8),
    to_signed(2, 8),
    to_signed(3, 8),
    to_signed(3, 8),
    to_signed(5, 8),
    to_signed(5, 8),
    to_signed(5, 8),
    to_signed(3, 8),
    to_signed(2, 8),
    to_signed(2, 8),
    to_signed(4, 8),
    to_signed(4, 8),
    to_signed(3, 8),
    to_signed(2, 8),
    to_signed(1, 8),
    to_signed(2, 8),
    to_signed(3, 8),
    to_signed(4, 8),
    to_signed(6, 8),
    to_signed(8, 8),
    to_signed(7, 8),
    to_signed(6, 8),
    to_signed(5, 8),
    to_signed(5, 8),
    to_signed(5, 8),
    to_signed(4, 8),
    to_signed(3, 8),
    to_signed(1, 8),
    to_signed(0, 8),
    to_signed(-2, 8),
    to_signed(-2, 8),
    to_signed(-2, 8),
    to_signed(-2, 8),
    to_signed(-1, 8),
    to_signed(0, 8),
    to_signed(1, 8),
    to_signed(2, 8),
    to_signed(1, 8),
    to_signed(1, 8),
    to_signed(1, 8),
    to_signed(2, 8),
    to_signed(3, 8),
    to_signed(4, 8),
    to_signed(4, 8),
    to_signed(6, 8),
    to_signed(6, 8),
    to_signed(6, 8),
    to_signed(6, 8),
    to_signed(6, 8),
    to_signed(4, 8),
    to_signed(2, 8),
    to_signed(1, 8),
    to_signed(0, 8),
    to_signed(1, 8),
    to_signed(3, 8),
    to_signed(6, 8),
    to_signed(7, 8),
    to_signed(6, 8),
    to_signed(5, 8),
    to_signed(4, 8),
    to_signed(4, 8),
    to_signed(4, 8),
    to_signed(3, 8),
    to_signed(3, 8),
    to_signed(4, 8),
    to_signed(6, 8),
    to_signed(7, 8),
    to_signed(7, 8),
    to_signed(5, 8),
    to_signed(4, 8),
    to_signed(3, 8),
    to_signed(1, 8),
    to_signed(-1, 8),
    to_signed(-2, 8),
    to_signed(-3, 8),
    to_signed(-2, 8),
    to_signed(0, 8),
    to_signed(1, 8),
    to_signed(3, 8),
    to_signed(4, 8),
    to_signed(4, 8),
    to_signed(5, 8),
    to_signed(5, 8),
    to_signed(4, 8),
    to_signed(3, 8),
    to_signed(3, 8),
    to_signed(4, 8),
    to_signed(5, 8),
    to_signed(6, 8),
    to_signed(6, 8),
    to_signed(6, 8),
    to_signed(5, 8),
    to_signed(3, 8),
    to_signed(2, 8),
    to_signed(1, 8),
    to_signed(0, 8),
    to_signed(-1, 8),
    to_signed(0, 8),
    to_signed(2, 8),
    to_signed(4, 8),
    to_signed(5, 8),
    to_signed(4, 8),
    to_signed(3, 8),
    to_signed(3, 8),
    to_signed(3, 8),
    to_signed(2, 8),
    to_signed(1, 8),
    to_signed(1, 8),
    to_signed(1, 8),
    to_signed(0, 8),
    to_signed(-1, 8),
    to_signed(-1, 8),
    to_signed(0, 8),
    to_signed(0, 8),
    to_signed(0, 8),
    to_signed(-1, 8),
    to_signed(-1, 8),
    to_signed(-2, 8),
    to_signed(-4, 8),
    to_signed(-4, 8),
    to_signed(-4, 8),
    to_signed(-3, 8),
    to_signed(-1, 8),
    to_signed(0, 8),
    to_signed(1, 8),
    to_signed(1, 8),
    to_signed(0, 8),
    to_signed(0, 8),
    to_signed(0, 8),
    to_signed(-1, 8),
    to_signed(-3, 8),
    to_signed(-5, 8),
    to_signed(-5, 8),
    to_signed(-4, 8),
    to_signed(-2, 8),
    to_signed(-1, 8),
    to_signed(0, 8),
    to_signed(0, 8),
    to_signed(-2, 8),
    to_signed(-4, 8),
    to_signed(-6, 8),
    to_signed(-6, 8),
    to_signed(-6, 8),
    to_signed(-5, 8),
    to_signed(-3, 8),
    to_signed(-3, 8),
    to_signed(-3, 8),
    to_signed(-4, 8),
    to_signed(-5, 8),
    to_signed(-5, 8),
    to_signed(-4, 8),
    to_signed(-5, 8),
    to_signed(-6, 8),
    to_signed(-7, 8),
    to_signed(-8, 8),
    to_signed(-7, 8),
    to_signed(-7, 8),
    to_signed(-6, 8),
    to_signed(-5, 8),
    to_signed(-5, 8),
    to_signed(-6, 8),
    to_signed(-7, 8),
    to_signed(-8, 8),
    to_signed(-8, 8),
    to_signed(-8, 8),
    to_signed(-7, 8),
    to_signed(-6, 8),
    to_signed(-6, 8),
    to_signed(-6, 8),
    to_signed(-6, 8),
    to_signed(-5, 8),
    to_signed(-4, 8),
    to_signed(-4, 8),
    to_signed(-5, 8),
    to_signed(-5, 8),
    to_signed(-6, 8),
    to_signed(-7, 8),
    to_signed(-7, 8),
    to_signed(-6, 8),
    to_signed(-5, 8),
    to_signed(-5, 8),
    to_signed(-4, 8),
    to_signed(-5, 8),
    to_signed(-6, 8),
    to_signed(-7, 8),
    to_signed(-7, 8),
    to_signed(-6, 8),
    to_signed(-4, 8),
    to_signed(-3, 8),
    to_signed(-4, 8),
    to_signed(-4, 8),
    to_signed(-5, 8),
    to_signed(-4, 8),
    to_signed(-4, 8),
    to_signed(-3, 8),
    to_signed(-1, 8),
    to_signed(0, 8),
    to_signed(-1, 8),
    to_signed(-3, 8),
    to_signed(-3, 8),
    to_signed(-4, 8),
    to_signed(-3, 8),
    to_signed(-3, 8),
    to_signed(-3, 8),
    to_signed(-2, 8),
    to_signed(-1, 8),
    to_signed(0, 8),
    to_signed(0, 8),
    to_signed(0, 8),
    to_signed(-1, 8),
    to_signed(-3, 8),
    to_signed(-4, 8),
    to_signed(-5, 8),
    to_signed(-4, 8),
    to_signed(-2, 8),
    to_signed(0, 8),
    to_signed(2, 8),
    to_signed(3, 8),
    to_signed(3, 8),
    to_signed(1, 8),
    to_signed(0, 8),
    to_signed(-2, 8),
    to_signed(-2, 8),
    to_signed(-1, 8),
    to_signed(0, 8),
    to_signed(-1, 8),
    to_signed(-2, 8),
    to_signed(-2, 8),
    to_signed(-1, 8),
    to_signed(1, 8),
    to_signed(1, 8),
    to_signed(0, 8),
    to_signed(-1, 8),
    to_signed(-2, 8),
    to_signed(-2, 8),
    to_signed(-1, 8),
    to_signed(1, 8),
    to_signed(4, 8),
    to_signed(6, 8),
    to_signed(7, 8),
    to_signed(7, 8),
    to_signed(7, 8),
    to_signed(6, 8),
    to_signed(5, 8),
    to_signed(4, 8),
    to_signed(4, 8),
    to_signed(3, 8),
    to_signed(2, 8),
    to_signed(2, 8),
    to_signed(2, 8),
    to_signed(3, 8),
    to_signed(4, 8),
    to_signed(5, 8),
    to_signed(3, 8),
    to_signed(2, 8),
    to_signed(1, 8),
    to_signed(1, 8),
    to_signed(3, 8),
    to_signed(4, 8),
    to_signed(6, 8),
    to_signed(7, 8),
    to_signed(7, 8),
    to_signed(6, 8),
    to_signed(5, 8),
    to_signed(4, 8),
    to_signed(4, 8),
    to_signed(3, 8),
    to_signed(2, 8),
    to_signed(1, 8),
    to_signed(-1, 8),
    to_signed(-3, 8),
    to_signed(-4, 8),
    to_signed(-4, 8),
    to_signed(-2, 8),
    to_signed(0, 8),
    to_signed(1, 8),
    to_signed(2, 8),
    to_signed(1, 8),
    to_signed(1, 8),
    to_signed(1, 8),
    to_signed(2, 8),
    to_signed(3, 8),
    to_signed(4, 8),
    to_signed(4, 8),
    to_signed(4, 8),
    to_signed(4, 8),
    to_signed(4, 8),
    to_signed(5, 8),
    to_signed(4, 8),
    to_signed(3, 8),
    to_signed(0, 8),
    to_signed(-2, 8),
    to_signed(-3, 8),
    to_signed(-3, 8),
    to_signed(-2, 8),
    to_signed(0, 8),
    to_signed(3, 8),
    to_signed(5, 8),
    to_signed(5, 8),
    to_signed(5, 8),
    to_signed(4, 8),
    to_signed(4, 8),
    to_signed(3, 8),
    to_signed(3, 8),
    to_signed(2, 8),
    to_signed(2, 8),
    to_signed(2, 8),
    to_signed(2, 8),
    to_signed(3, 8),
    to_signed(3, 8),
    to_signed(3, 8),
    to_signed(1, 8),
    to_signed(-2, 8),
    to_signed(-5, 8),
    to_signed(-8, 8),
    to_signed(-9, 8),
    to_signed(-8, 8),
    to_signed(-6, 8),
    to_signed(-2, 8),
    to_signed(0, 8),
    to_signed(2, 8),
    to_signed(2, 8),
    to_signed(1, 8),
    to_signed(-1, 8),
    to_signed(-2, 8),
    to_signed(-2, 8),
    to_signed(-2, 8),
    to_signed(-2, 8),
    to_signed(-1, 8),
    to_signed(0, 8),
    to_signed(0, 8),
    to_signed(0, 8),
    to_signed(0, 8),
    to_signed(-1, 8),
    to_signed(-3, 8),
    to_signed(-5, 8),
    to_signed(-6, 8),
    to_signed(-5, 8),
    to_signed(-3, 8),
    to_signed(1, 8),
    to_signed(4, 8),
    to_signed(5, 8),
    to_signed(5, 8),
    to_signed(4, 8),
    to_signed(4, 8),
    to_signed(3, 8),
    to_signed(4, 8),
    to_signed(4, 8),
    to_signed(5, 8),
    to_signed(4, 8),
    to_signed(3, 8),
    to_signed(2, 8),
    to_signed(2, 8),
    to_signed(3, 8),
    to_signed(4, 8),
    to_signed(4, 8),
    to_signed(4, 8),
    to_signed(3, 8),
    to_signed(1, 8),
    to_signed(-1, 8),
    to_signed(-2, 8),
    to_signed(-1, 8),
    to_signed(1, 8),
    to_signed(2, 8),
    to_signed(3, 8),
    to_signed(3, 8),
    to_signed(3, 8),
    to_signed(3, 8),
    to_signed(3, 8),
    to_signed(2, 8),
    to_signed(0, 8),
    to_signed(-2, 8),
    to_signed(-4, 8),
    to_signed(-6, 8),
    to_signed(-8, 8),
    to_signed(-7, 8),
    to_signed(-6, 8),
    to_signed(-3, 8),
    to_signed(-1, 8),
    to_signed(-1, 8),
    to_signed(-1, 8),
    to_signed(-1, 8),
    to_signed(-2, 8),
    to_signed(-4, 8),
    to_signed(-5, 8),
    to_signed(-5, 8),
    to_signed(-5, 8),
    to_signed(-4, 8),
    to_signed(-2, 8),
    to_signed(0, 8),
    to_signed(2, 8),
    to_signed(2, 8),
    to_signed(0, 8),
    to_signed(-4, 8),
    to_signed(-7, 8),
    to_signed(-10, 8),
    to_signed(-10, 8),
    to_signed(-8, 8),
    to_signed(-4, 8),
    to_signed(-1, 8),
    to_signed(1, 8),
    to_signed(1, 8),
    to_signed(0, 8),
    to_signed(-1, 8),
    to_signed(-3, 8),
    to_signed(-4, 8),
    to_signed(-5, 8),
    to_signed(-4, 8),
    to_signed(-3, 8),
    to_signed(0, 8),
    to_signed(2, 8),
    to_signed(5, 8),
    to_signed(6, 8),
    to_signed(6, 8),
    to_signed(5, 8),
    to_signed(4, 8),
    to_signed(4, 8),
    to_signed(3, 8),
    to_signed(3, 8),
    to_signed(3, 8),
    to_signed(4, 8),
    to_signed(6, 8),
    to_signed(7, 8),
    to_signed(7, 8),
    to_signed(7, 8),
    to_signed(6, 8),
    to_signed(6, 8),
    to_signed(6, 8),
    to_signed(5, 8),
    to_signed(3, 8),
    to_signed(1, 8),
    to_signed(0, 8),
    to_signed(2, 8),
    to_signed(4, 8),
    to_signed(6, 8),
    to_signed(7, 8),
    to_signed(7, 8),
    to_signed(6, 8),
    to_signed(4, 8),
    to_signed(3, 8),
    to_signed(1, 8),
    to_signed(0, 8),
    to_signed(0, 8),
    to_signed(0, 8),
    to_signed(0, 8),
    to_signed(0, 8),
    to_signed(0, 8),
    to_signed(0, 8),
    to_signed(1, 8),
    to_signed(1, 8),
    to_signed(-1, 8),
    to_signed(-3, 8),
    to_signed(-5, 8),
    to_signed(-4, 8),
    to_signed(-3, 8),
    to_signed(0, 8),
    to_signed(3, 8),
    to_signed(6, 8),
    to_signed(8, 8),
    to_signed(9, 8),
    to_signed(8, 8),
    to_signed(6, 8),
    to_signed(3, 8),
    to_signed(1, 8),
    to_signed(1, 8),
    to_signed(1, 8),
    to_signed(1, 8),
    to_signed(3, 8),
    to_signed(5, 8),
    to_signed(7, 8),
    to_signed(8, 8),
    to_signed(6, 8),
    to_signed(4, 8),
    to_signed(2, 8),
    to_signed(0, 8),
    to_signed(-1, 8),
    to_signed(0, 8),
    to_signed(3, 8),
    to_signed(6, 8),
    to_signed(9, 8),
    to_signed(10, 8),
    to_signed(10, 8),
    to_signed(10, 8),
    to_signed(8, 8),
    to_signed(5, 8),
    to_signed(1, 8),
    to_signed(-3, 8),
    to_signed(-4, 8),
    to_signed(-4, 8),
    to_signed(-4, 8),
    to_signed(-4, 8),
    to_signed(-4, 8),
    to_signed(-4, 8),
    to_signed(-3, 8),
    to_signed(-4, 8),
    to_signed(-7, 8),
    to_signed(-9, 8),
    to_signed(-9, 8),
    to_signed(-7, 8),
    to_signed(-5, 8),
    to_signed(-4, 8),
    to_signed(-4, 8),
    to_signed(-3, 8),
    to_signed(-1, 8),
    to_signed(0, 8),
    to_signed(-2, 8),
    to_signed(-5, 8),
    to_signed(-8, 8),
    to_signed(-9, 8),
    to_signed(-11, 8),
    to_signed(-11, 8),
    to_signed(-10, 8),
    to_signed(-8, 8),
    to_signed(-6, 8),
    to_signed(-6, 8),
    to_signed(-6, 8),
    to_signed(-7, 8),
    to_signed(-7, 8),
    to_signed(-7, 8),
    to_signed(-6, 8),
    to_signed(-4, 8),
    to_signed(-3, 8),
    to_signed(-2, 8),
    to_signed(0, 8),
    to_signed(3, 8),
    to_signed(6, 8),
    to_signed(7, 8),
    to_signed(6, 8),
    to_signed(3, 8),
    to_signed(0, 8),
    to_signed(-3, 8),
    to_signed(-6, 8),
    to_signed(-6, 8),
    to_signed(-4, 8),
    to_signed(-2, 8),
    to_signed(1, 8),
    to_signed(2, 8),
    to_signed(2, 8),
    to_signed(2, 8),
    to_signed(1, 8),
    to_signed(0, 8),
    to_signed(-1, 8),
    to_signed(-1, 8),
    to_signed(-1, 8),
    to_signed(-1, 8),
    to_signed(-1, 8),
    to_signed(-1, 8),
    to_signed(0, 8),
    to_signed(2, 8),
    to_signed(3, 8),
    to_signed(2, 8),
    to_signed(-1, 8),
    to_signed(-5, 8),
    to_signed(-8, 8),
    to_signed(-10, 8),
    to_signed(-11, 8),
    to_signed(-9, 8),
    to_signed(-8, 8),
    to_signed(-6, 8),
    to_signed(-5, 8),
    to_signed(-4, 8),
    to_signed(-4, 8),
    to_signed(-4, 8),
    to_signed(-5, 8),
    to_signed(-6, 8),
    to_signed(-7, 8),
    to_signed(-7, 8),
    to_signed(-6, 8),
    to_signed(-4, 8),
    to_signed(-1, 8),
    to_signed(1, 8),
    to_signed(1, 8),
    to_signed(0, 8),
    to_signed(-1, 8),
    to_signed(-3, 8),
    to_signed(-5, 8),
    to_signed(-6, 8),
    to_signed(-6, 8),
    to_signed(-4, 8),
    to_signed(-2, 8),
    to_signed(-1, 8),
    to_signed(0, 8),
    to_signed(1, 8),
    to_signed(2, 8),
    to_signed(3, 8),
    to_signed(2, 8),
    to_signed(1, 8),
    to_signed(-1, 8),
    to_signed(-2, 8),
    to_signed(-2, 8),
    to_signed(-1, 8),
    to_signed(1, 8),
    to_signed(2, 8),
    to_signed(4, 8),
    to_signed(4, 8),
    to_signed(2, 8),
    to_signed(0, 8),
    to_signed(-3, 8),
    to_signed(-4, 8),
    to_signed(-5, 8),
    to_signed(-6, 8),
    to_signed(-6, 8),
    to_signed(-4, 8),
    to_signed(-2, 8),
    to_signed(0, 8),
    to_signed(-1, 8),
    to_signed(-3, 8),
    to_signed(-4, 8),
    to_signed(-5, 8),
    to_signed(-6, 8),
    to_signed(-7, 8),
    to_signed(-7, 8),
    to_signed(-6, 8),
    to_signed(-4, 8),
    to_signed(-2, 8),
    to_signed(-1, 8),
    to_signed(-1, 8),
    to_signed(-1, 8),
    to_signed(-2, 8),
    to_signed(-4, 8),
    to_signed(-6, 8),
    to_signed(-6, 8),
    to_signed(-7, 8),
    to_signed(-7, 8),
    to_signed(-6, 8),
    to_signed(-6, 8),
    to_signed(-5, 8),
    to_signed(-3, 8),
    to_signed(-2, 8),
    to_signed(-2, 8),
    to_signed(-3, 8),
    to_signed(-4, 8),
    to_signed(-5, 8),
    to_signed(-6, 8),
    to_signed(-6, 8),
    to_signed(-4, 8),
    to_signed(-2, 8),
    to_signed(-1, 8),
    to_signed(-1, 8),
    to_signed(0, 8),
    to_signed(0, 8),
    to_signed(-1, 8),
    to_signed(-3, 8),
    to_signed(-6, 8),
    to_signed(-8, 8),
    to_signed(-9, 8),
    to_signed(-10, 8),
    to_signed(-10, 8),
    to_signed(-9, 8),
    to_signed(-7, 8),
    to_signed(-5, 8),
    to_signed(-3, 8),
    to_signed(-3, 8),
    to_signed(-3, 8),
    to_signed(-4, 8),
    to_signed(-5, 8),
    to_signed(-5, 8),
    to_signed(-5, 8),
    to_signed(-3, 8),
    to_signed(-1, 8),
    to_signed(1, 8),
    to_signed(2, 8),
    to_signed(2, 8),
    to_signed(1, 8),
    to_signed(-1, 8),
    to_signed(-3, 8),
    to_signed(-6, 8),
    to_signed(-9, 8),
    to_signed(-11, 8),
    to_signed(-10, 8),
    to_signed(-8, 8),
    to_signed(-4, 8),
    to_signed(-2, 8),
    to_signed(-1, 8),
    to_signed(0, 8),
    to_signed(0, 8),
    to_signed(-2, 8),
    to_signed(-3, 8),
    to_signed(-3, 8),
    to_signed(-1, 8),
    to_signed(2, 8),
    to_signed(4, 8),
    to_signed(6, 8),
    to_signed(7, 8),
    to_signed(7, 8),
    to_signed(6, 8),
    to_signed(3, 8),
    to_signed(0, 8),
    to_signed(-1, 8),
    to_signed(-2, 8),
    to_signed(-3, 8),
    to_signed(-2, 8),
    to_signed(0, 8),
    to_signed(3, 8),
    to_signed(6, 8),
    to_signed(8, 8),
    to_signed(8, 8),
    to_signed(7, 8),
    to_signed(5, 8),
    to_signed(4, 8),
    to_signed(4, 8),
    to_signed(6, 8),
    to_signed(7, 8),
    to_signed(8, 8),
    to_signed(8, 8),
    to_signed(8, 8),
    to_signed(7, 8),
    to_signed(6, 8),
    to_signed(3, 8),
    to_signed(0, 8),
    to_signed(-3, 8),
    to_signed(-5, 8),
    to_signed(-6, 8),
    to_signed(-6, 8),
    to_signed(-6, 8),
    to_signed(-4, 8),
    to_signed(-1, 8),
    to_signed(0, 8),
    to_signed(0, 8),
    to_signed(-1, 8),
    to_signed(-1, 8),
    to_signed(-2, 8),
    to_signed(-3, 8),
    to_signed(-4, 8),
    to_signed(-3, 8),
    to_signed(-2, 8),
    to_signed(-1, 8),
    to_signed(-1, 8),
    to_signed(-2, 8),
    to_signed(-3, 8),
    to_signed(-3, 8),
    to_signed(-4, 8),
    to_signed(-4, 8),
    to_signed(-5, 8),
    to_signed(-6, 8),
    to_signed(-7, 8),
    to_signed(-5, 8),
    to_signed(-3, 8),
    to_signed(-1, 8),
    to_signed(0, 8),
    to_signed(2, 8),
    to_signed(4, 8),
    to_signed(5, 8),
    to_signed(5, 8),
    to_signed(5, 8),
    to_signed(4, 8),
    to_signed(2, 8),
    to_signed(0, 8),
    to_signed(1, 8),
    to_signed(3, 8),
    to_signed(5, 8),
    to_signed(6, 8),
    to_signed(6, 8),
    to_signed(4, 8),
    to_signed(3, 8),
    to_signed(1, 8),
    to_signed(-1, 8),
    to_signed(-2, 8),
    to_signed(-2, 8),
    to_signed(-1, 8),
    to_signed(2, 8),
    to_signed(4, 8),
    to_signed(7, 8),
    to_signed(9, 8),
    to_signed(9, 8),
    to_signed(7, 8),
    to_signed(5, 8),
    to_signed(1, 8),
    to_signed(-2, 8),
    to_signed(-4, 8),
    to_signed(-3, 8),
    to_signed(-2, 8),
    to_signed(0, 8),
    to_signed(2, 8),
    to_signed(3, 8),
    to_signed(4, 8),
    to_signed(2, 8),
    to_signed(0, 8),
    to_signed(-4, 8),
    to_signed(-7, 8),
    to_signed(-8, 8),
    to_signed(-8, 8),
    to_signed(-6, 8),
    to_signed(-4, 8),
    to_signed(-2, 8),
    to_signed(0, 8),
    to_signed(1, 8),
    to_signed(1, 8),
    to_signed(0, 8),
    to_signed(-2, 8),
    to_signed(-5, 8),
    to_signed(-6, 8),
    to_signed(-6, 8),
    to_signed(-5, 8),
    to_signed(-3, 8),
    to_signed(-1, 8),
    to_signed(1, 8),
    to_signed(2, 8),
    to_signed(1, 8),
    to_signed(-1, 8),
    to_signed(-3, 8),
    to_signed(-6, 8),
    to_signed(-8, 8),
    to_signed(-9, 8),
    to_signed(-7, 8),
    to_signed(-4, 8),
    to_signed(-1, 8),
    to_signed(1, 8),
    to_signed(2, 8),
    to_signed(2, 8),
    to_signed(2, 8),
    to_signed(2, 8),
    to_signed(1, 8),
    to_signed(0, 8),
    to_signed(0, 8),
    to_signed(1, 8),
    to_signed(2, 8),
    to_signed(3, 8),
    to_signed(3, 8),
    to_signed(2, 8),
    to_signed(2, 8),
    to_signed(2, 8),
    to_signed(1, 8),
    to_signed(-1, 8),
    to_signed(-3, 8),
    to_signed(-4, 8),
    to_signed(-4, 8),
    to_signed(-2, 8),
    to_signed(-1, 8),
    to_signed(1, 8),
    to_signed(3, 8),
    to_signed(3, 8),
    to_signed(3, 8),
    to_signed(3, 8),
    to_signed(2, 8),
    to_signed(2, 8),
    to_signed(1, 8),
    to_signed(0, 8),
    to_signed(-1, 8),
    to_signed(0, 8),
    to_signed(1, 8),
    to_signed(3, 8),
    to_signed(3, 8),
    to_signed(2, 8),
    to_signed(-1, 8),
    to_signed(-5, 8),
    to_signed(-8, 8),
    to_signed(-9, 8),
    to_signed(-9, 8),
    to_signed(-7, 8),
    to_signed(-5, 8),
    to_signed(-3, 8),
    to_signed(-1, 8),
    to_signed(1, 8),
    to_signed(2, 8),
    to_signed(3, 8),
    to_signed(2, 8),
    to_signed(0, 8),
    to_signed(-1, 8),
    to_signed(-2, 8),
    to_signed(-2, 8),
    to_signed(-2, 8),
    to_signed(-2, 8),
    to_signed(-2, 8),
    to_signed(-2, 8),
    to_signed(-2, 8),
    to_signed(-3, 8),
    to_signed(-4, 8),
    to_signed(-7, 8),
    to_signed(-10, 8),
    to_signed(-12, 8),
    to_signed(-10, 8),
    to_signed(-7, 8),
    to_signed(-4, 8),
    to_signed(-1, 8),
    to_signed(1, 8),
    to_signed(3, 8),
    to_signed(4, 8),
    to_signed(4, 8),
    to_signed(2, 8),
    to_signed(0, 8),
    to_signed(-2, 8),
    to_signed(-3, 8),
    to_signed(-5, 8),
    to_signed(-5, 8),
    to_signed(-4, 8),
    to_signed(-2, 8),
    to_signed(-1, 8),
    to_signed(-1, 8),
    to_signed(-3, 8),
    to_signed(-5, 8),
    to_signed(-6, 8),
    to_signed(-5, 8),
    to_signed(-2, 8),
    to_signed(2, 8),
    to_signed(4, 8),
    to_signed(6, 8),
    to_signed(7, 8),
    to_signed(8, 8),
    to_signed(8, 8),
    to_signed(8, 8),
    to_signed(7, 8),
    to_signed(5, 8),
    to_signed(3, 8),
    to_signed(1, 8),
    to_signed(0, 8),
    to_signed(0, 8),
    to_signed(0, 8),
    to_signed(2, 8),
    to_signed(2, 8),
    to_signed(1, 8),
    to_signed(-2, 8),
    to_signed(-4, 8),
    to_signed(-5, 8),
    to_signed(-4, 8),
    to_signed(-3, 8),
    to_signed(-1, 8),
    to_signed(0, 8),
    to_signed(1, 8),
    to_signed(1, 8),
    to_signed(2, 8),
    to_signed(2, 8),
    to_signed(2, 8),
    to_signed(1, 8),
    to_signed(-1, 8),
    to_signed(-5, 8),
    to_signed(-8, 8),
    to_signed(-9, 8),
    to_signed(-8, 8),
    to_signed(-6, 8),
    to_signed(-3, 8),
    to_signed(-2, 8),
    to_signed(-3, 8),
    to_signed(-4, 8),
    to_signed(-6, 8),
    to_signed(-7, 8),
    to_signed(-8, 8),
    to_signed(-7, 8),
    to_signed(-5, 8),
    to_signed(-3, 8),
    to_signed(-2, 8),
    to_signed(-1, 8),
    to_signed(0, 8),
    to_signed(1, 8),
    to_signed(1, 8),
    to_signed(1, 8),
    to_signed(0, 8),
    to_signed(-1, 8),
    to_signed(-2, 8),
    to_signed(-4, 8),
    to_signed(-4, 8),
    to_signed(-3, 8),
    to_signed(-1, 8),
    to_signed(2, 8),
    to_signed(3, 8),
    to_signed(4, 8),
    to_signed(4, 8),
    to_signed(4, 8),
    to_signed(2, 8),
    to_signed(1, 8),
    to_signed(2, 8),
    to_signed(2, 8),
    to_signed(4, 8),
    to_signed(5, 8),
    to_signed(7, 8),
    to_signed(10, 8),
    to_signed(12, 8),
    to_signed(12, 8),
    to_signed(10, 8),
    to_signed(8, 8),
    to_signed(6, 8),
    to_signed(4, 8),
    to_signed(4, 8),
    to_signed(4, 8),
    to_signed(6, 8),
    to_signed(9, 8),
    to_signed(11, 8),
    to_signed(11, 8),
    to_signed(8, 8),
    to_signed(4, 8),
    to_signed(2, 8),
    to_signed(0, 8),
    to_signed(0, 8),
    to_signed(-1, 8),
    to_signed(1, 8),
    to_signed(3, 8),
    to_signed(5, 8),
    to_signed(6, 8),
    to_signed(6, 8),
    to_signed(5, 8),
    to_signed(4, 8),
    to_signed(1, 8),
    to_signed(-1, 8),
    to_signed(-4, 8),
    to_signed(-4, 8),
    to_signed(-3, 8),
    to_signed(-2, 8),
    to_signed(-1, 8),
    to_signed(0, 8),
    to_signed(1, 8),
    to_signed(0, 8),
    to_signed(-2, 8),
    to_signed(-5, 8),
    to_signed(-8, 8),
    to_signed(-10, 8),
    to_signed(-10, 8),
    to_signed(-7, 8),
    to_signed(-4, 8),
    to_signed(0, 8),
    to_signed(4, 8),
    to_signed(6, 8),
    to_signed(5, 8),
    to_signed(3, 8),
    to_signed(1, 8),
    to_signed(0, 8),
    to_signed(-1, 8),
    to_signed(-1, 8),
    to_signed(-1, 8),
    to_signed(1, 8),
    to_signed(4, 8),
    to_signed(6, 8),
    to_signed(7, 8),
    to_signed(7, 8),
    to_signed(5, 8),
    to_signed(3, 8),
    to_signed(2, 8),
    to_signed(2, 8),
    to_signed(3, 8),
    to_signed(5, 8),
    to_signed(6, 8),
    to_signed(8, 8),
    to_signed(10, 8),
    to_signed(12, 8),
    to_signed(12, 8),
    to_signed(11, 8),
    to_signed(10, 8),
    to_signed(7, 8),
    to_signed(4, 8),
    to_signed(1, 8),
    to_signed(0, 8),
    to_signed(1, 8),
    to_signed(1, 8),
    to_signed(1, 8),
    to_signed(0, 8),
    to_signed(-2, 8),
    to_signed(-4, 8),
    to_signed(-5, 8),
    to_signed(-5, 8),
    to_signed(-5, 8),
    to_signed(-5, 8),
    to_signed(-5, 8),
    to_signed(-5, 8),
    to_signed(-2, 8),
    to_signed(1, 8),
    to_signed(5, 8),
    to_signed(6, 8),
    to_signed(5, 8),
    to_signed(3, 8),
    to_signed(0, 8),
    to_signed(-4, 8),
    to_signed(-6, 8),
    to_signed(-6, 8),
    to_signed(-3, 8),
    to_signed(0, 8),
    to_signed(2, 8),
    to_signed(0, 8),
    to_signed(-1, 8),
    to_signed(-2, 8),
    to_signed(-1, 8),
    to_signed(0, 8),
    to_signed(1, 8),
    to_signed(1, 8),
    to_signed(1, 8),
    to_signed(0, 8),
    to_signed(2, 8),
    to_signed(5, 8),
    to_signed(9, 8),
    to_signed(13, 8),
    to_signed(14, 8),
    to_signed(13, 8),
    to_signed(8, 8),
    to_signed(2, 8),
    to_signed(-2, 8),
    to_signed(-4, 8),
    to_signed(-2, 8),
    to_signed(1, 8),
    to_signed(5, 8),
    to_signed(7, 8),
    to_signed(7, 8),
    to_signed(6, 8),
    to_signed(4, 8),
    to_signed(3, 8),
    to_signed(2, 8),
    to_signed(2, 8),
    to_signed(1, 8),
    to_signed(1, 8),
    to_signed(3, 8),
    to_signed(5, 8),
    to_signed(9, 8),
    to_signed(13, 8),
    to_signed(15, 8),
    to_signed(13, 8),
    to_signed(8, 8),
    to_signed(1, 8),
    to_signed(-4, 8),
    to_signed(-6, 8),
    to_signed(-5, 8),
    to_signed(-2, 8),
    to_signed(0, 8),
    to_signed(2, 8),
    to_signed(3, 8),
    to_signed(3, 8),
    to_signed(3, 8),
    to_signed(3, 8),
    to_signed(2, 8),
    to_signed(0, 8),
    to_signed(-3, 8),
    to_signed(-4, 8),
    to_signed(-5, 8),
    to_signed(-2, 8),
    to_signed(2, 8),
    to_signed(5, 8),
    to_signed(6, 8),
    to_signed(4, 8),
    to_signed(0, 8),
    to_signed(-4, 8),
    to_signed(-8, 8),
    to_signed(-9, 8),
    to_signed(-8, 8),
    to_signed(-5, 8),
    to_signed(-3, 8),
    to_signed(-1, 8),
    to_signed(-1, 8),
    to_signed(-1, 8),
    to_signed(-2, 8),
    to_signed(-3, 8),
    to_signed(-5, 8),
    to_signed(-8, 8),
    to_signed(-10, 8),
    to_signed(-9, 8),
    to_signed(-7, 8),
    to_signed(-4, 8),
    to_signed(-1, 8),
    to_signed(1, 8),
    to_signed(0, 8),
    to_signed(-3, 8),
    to_signed(-6, 8),
    to_signed(-8, 8),
    to_signed(-8, 8),
    to_signed(-7, 8),
    to_signed(-6, 8),
    to_signed(-5, 8),
    to_signed(-5, 8),
    to_signed(-7, 8),
    to_signed(-9, 8),
    to_signed(-7, 8),
    to_signed(-5, 8),
    to_signed(-4, 8),
    to_signed(-7, 8),
    to_signed(-12, 8),
    to_signed(-15, 8),
    to_signed(-15, 8),
    to_signed(-12, 8),
    to_signed(-8, 8),
    to_signed(-3, 8),
    to_signed(1, 8),
    to_signed(3, 8),
    to_signed(3, 8),
    to_signed(1, 8),
    to_signed(-1, 8),
    to_signed(-3, 8),
    to_signed(-4, 8),
    to_signed(-4, 8),
    to_signed(-4, 8),
    to_signed(-4, 8),
    to_signed(-4, 8),
    to_signed(-4, 8),
    to_signed(-3, 8),
    to_signed(-1, 8),
    to_signed(1, 8),
    to_signed(1, 8),
    to_signed(-1, 8),
    to_signed(-4, 8),
    to_signed(-7, 8),
    to_signed(-8, 8),
    to_signed(-6, 8),
    to_signed(-2, 8),
    to_signed(2, 8),
    to_signed(3, 8),
    to_signed(3, 8),
    to_signed(1, 8),
    to_signed(-1, 8),
    to_signed(-3, 8),
    to_signed(-5, 8),
    to_signed(-7, 8),
    to_signed(-9, 8),
    to_signed(-11, 8),
    to_signed(-11, 8),
    to_signed(-9, 8),
    to_signed(-7, 8),
    to_signed(-6, 8),
    to_signed(-4, 8),
    to_signed(-5, 8),
    to_signed(-6, 8),
    to_signed(-8, 8),
    to_signed(-10, 8),
    to_signed(-10, 8),
    to_signed(-8, 8),
    to_signed(-5, 8),
    to_signed(-3, 8),
    to_signed(-1, 8),
    to_signed(1, 8),
    to_signed(0, 8),
    to_signed(-2, 8),
    to_signed(-4, 8),
    to_signed(-5, 8),
    to_signed(-6, 8),
    to_signed(-6, 8),
    to_signed(-7, 8),
    to_signed(-6, 8),
    to_signed(-5, 8),
    to_signed(-3, 8),
    to_signed(-2, 8),
    to_signed(-1, 8),
    to_signed(-1, 8),
    to_signed(-1, 8),
    to_signed(-3, 8),
    to_signed(-4, 8),
    to_signed(-3, 8),
    to_signed(-1, 8),
    to_signed(0, 8),
    to_signed(2, 8),
    to_signed(4, 8),
    to_signed(7, 8),
    to_signed(9, 8),
    to_signed(7, 8),
    to_signed(4, 8),
    to_signed(1, 8),
    to_signed(-3, 8),
    to_signed(-6, 8),
    to_signed(-7, 8),
    to_signed(-7, 8),
    to_signed(-5, 8),
    to_signed(-4, 8),
    to_signed(-2, 8),
    to_signed(-2, 8),
    to_signed(-3, 8),
    to_signed(-6, 8),
    to_signed(-8, 8),
    to_signed(-8, 8),
    to_signed(-8, 8),
    to_signed(-8, 8),
    to_signed(-7, 8),
    to_signed(-5, 8),
    to_signed(-4, 8),
    to_signed(-2, 8),
    to_signed(-2, 8),
    to_signed(-3, 8),
    to_signed(-5, 8),
    to_signed(-6, 8),
    to_signed(-8, 8),
    to_signed(-9, 8),
    to_signed(-10, 8),
    to_signed(-11, 8),
    to_signed(-10, 8),
    to_signed(-8, 8),
    to_signed(-7, 8),
    to_signed(-5, 8),
    to_signed(-2, 8),
    to_signed(0, 8),
    to_signed(-1, 8),
    to_signed(-2, 8),
    to_signed(-3, 8),
    to_signed(-2, 8),
    to_signed(-1, 8),
    to_signed(0, 8),
    to_signed(2, 8),
    to_signed(3, 8),
    to_signed(4, 8),
    to_signed(3, 8),
    to_signed(2, 8),
    to_signed(1, 8),
    to_signed(1, 8),
    to_signed(2, 8),
    to_signed(2, 8),
    to_signed(2, 8),
    to_signed(1, 8),
    to_signed(0, 8),
    to_signed(1, 8),
    to_signed(2, 8),
    to_signed(4, 8),
    to_signed(5, 8),
    to_signed(5, 8),
    to_signed(4, 8),
    to_signed(2, 8),
    to_signed(0, 8),
    to_signed(-1, 8),
    to_signed(-1, 8),
    to_signed(1, 8),
    to_signed(3, 8),
    to_signed(4, 8),
    to_signed(5, 8),
    to_signed(5, 8),
    to_signed(5, 8),
    to_signed(3, 8),
    to_signed(2, 8),
    to_signed(0, 8),
    to_signed(-2, 8),
    to_signed(-3, 8),
    to_signed(-2, 8),
    to_signed(-1, 8),
    to_signed(1, 8),
    to_signed(3, 8),
    to_signed(3, 8),
    to_signed(2, 8),
    to_signed(-1, 8),
    to_signed(-3, 8),
    to_signed(-4, 8),
    to_signed(-4, 8),
    to_signed(-3, 8),
    to_signed(0, 8),
    to_signed(2, 8),
    to_signed(3, 8),
    to_signed(2, 8),
    to_signed(1, 8),
    to_signed(0, 8),
    to_signed(1, 8),
    to_signed(2, 8),
    to_signed(1, 8),
    to_signed(0, 8),
    to_signed(-1, 8),
    to_signed(-1, 8),
    to_signed(0, 8),
    to_signed(2, 8),
    to_signed(5, 8),
    to_signed(7, 8),
    to_signed(8, 8),
    to_signed(8, 8),
    to_signed(8, 8),
    to_signed(6, 8),
    to_signed(5, 8),
    to_signed(4, 8),
    to_signed(5, 8),
    to_signed(8, 8),
    to_signed(10, 8),
    to_signed(11, 8),
    to_signed(12, 8),
    to_signed(12, 8),
    to_signed(11, 8),
    to_signed(9, 8),
    to_signed(6, 8),
    to_signed(3, 8),
    to_signed(1, 8),
    to_signed(1, 8),
    to_signed(2, 8),
    to_signed(4, 8),
    to_signed(6, 8),
    to_signed(6, 8),
    to_signed(5, 8),
    to_signed(4, 8),
    to_signed(3, 8),
    to_signed(3, 8),
    to_signed(3, 8),
    to_signed(4, 8),
    to_signed(5, 8),
    to_signed(5, 8),
    to_signed(6, 8),
    to_signed(6, 8),
    to_signed(5, 8),
    to_signed(4, 8),
    to_signed(3, 8),
    to_signed(1, 8),
    to_signed(-1, 8),
    to_signed(-3, 8),
    to_signed(-5, 8),
    to_signed(-4, 8),
    to_signed(-2, 8),
    to_signed(-1, 8),
    to_signed(-1, 8),
    to_signed(-1, 8),
    to_signed(0, 8),
    to_signed(1, 8),
    to_signed(2, 8),
    to_signed(2, 8),
    to_signed(3, 8),
    to_signed(3, 8),
    to_signed(2, 8),
    to_signed(2, 8),
    to_signed(4, 8),
    to_signed(6, 8),
    to_signed(8, 8),
    to_signed(7, 8),
    to_signed(4, 8),
    to_signed(2, 8),
    to_signed(1, 8),
    to_signed(0, 8),
    to_signed(0, 8),
    to_signed(-1, 8),
    to_signed(0, 8),
    to_signed(1, 8),
    to_signed(2, 8),
    to_signed(3, 8),
    to_signed(4, 8),
    to_signed(5, 8),
    to_signed(5, 8),
    to_signed(4, 8),
    to_signed(1, 8),
    to_signed(-1, 8),
    to_signed(-1, 8),
    to_signed(1, 8),
    to_signed(3, 8),
    to_signed(4, 8),
    to_signed(5, 8),
    to_signed(4, 8),
    to_signed(3, 8),
    to_signed(-1, 8),
    to_signed(-5, 8),
    to_signed(-9, 8),
    to_signed(-10, 8),
    to_signed(-9, 8),
    to_signed(-7, 8),
    to_signed(-5, 8),
    to_signed(-5, 8),
    to_signed(-4, 8),
    to_signed(-3, 8),
    to_signed(-3, 8),
    to_signed(-3, 8),
    to_signed(-4, 8),
    to_signed(-5, 8),
    to_signed(-6, 8),
    to_signed(-7, 8),
    to_signed(-6, 8),
    to_signed(-5, 8),
    to_signed(-3, 8),
    to_signed(-2, 8),
    to_signed(-2, 8),
    to_signed(-3, 8),
    to_signed(-4, 8),
    to_signed(-5, 8),
    to_signed(-6, 8),
    to_signed(-7, 8),
    to_signed(-6, 8),
    to_signed(-5, 8),
    to_signed(-5, 8),
    to_signed(-4, 8),
    to_signed(-3, 8),
    to_signed(-3, 8),
    to_signed(-3, 8),
    to_signed(-4, 8),
    to_signed(-4, 8),
    to_signed(-4, 8),
    to_signed(-5, 8),
    to_signed(-6, 8),
    to_signed(-4, 8),
    to_signed(-2, 8),
    to_signed(0, 8),
    to_signed(0, 8),
    to_signed(1, 8),
    to_signed(1, 8),
    to_signed(0, 8),
    to_signed(-3, 8),
    to_signed(-5, 8),
    to_signed(-8, 8),
    to_signed(-9, 8),
    to_signed(-10, 8),
    to_signed(-9, 8),
    to_signed(-6, 8),
    to_signed(-3, 8),
    to_signed(-2, 8),
    to_signed(-2, 8),
    to_signed(-3, 8),
    to_signed(-5, 8),
    to_signed(-6, 8),
    to_signed(-7, 8),
    to_signed(-8, 8),
    to_signed(-8, 8),
    to_signed(-6, 8),
    to_signed(-2, 8),
    to_signed(0, 8),
    to_signed(1, 8),
    to_signed(-1, 8),
    to_signed(-4, 8),
    to_signed(-7, 8),
    to_signed(-10, 8),
    to_signed(-13, 8),
    to_signed(-15, 8),
    to_signed(-13, 8),
    to_signed(-11, 8),
    to_signed(-8, 8),
    to_signed(-5, 8),
    to_signed(-2, 8),
    to_signed(0, 8),
    to_signed(-1, 8),
    to_signed(-2, 8),
    to_signed(-4, 8),
    to_signed(-5, 8),
    to_signed(-4, 8),
    to_signed(-2, 8),
    to_signed(0, 8),
    to_signed(3, 8),
    to_signed(4, 8),
    to_signed(5, 8),
    to_signed(6, 8),
    to_signed(5, 8),
    to_signed(3, 8),
    to_signed(0, 8),
    to_signed(-3, 8),
    to_signed(-5, 8),
    to_signed(-4, 8),
    to_signed(-3, 8),
    to_signed(-2, 8),
    to_signed(1, 8),
    to_signed(4, 8),
    to_signed(5, 8),
    to_signed(5, 8),
    to_signed(3, 8),
    to_signed(2, 8),
    to_signed(2, 8),
    to_signed(3, 8),
    to_signed(4, 8),
    to_signed(5, 8),
    to_signed(7, 8),
    to_signed(10, 8),
    to_signed(10, 8),
    to_signed(9, 8),
    to_signed(5, 8),
    to_signed(1, 8),
    to_signed(-3, 8),
    to_signed(-6, 8),
    to_signed(-7, 8),
    to_signed(-5, 8),
    to_signed(-2, 8),
    to_signed(0, 8),
    to_signed(1, 8),
    to_signed(1, 8),
    to_signed(2, 8),
    to_signed(3, 8),
    to_signed(2, 8),
    to_signed(1, 8),
    to_signed(1, 8),
    to_signed(1, 8),
    to_signed(1, 8),
    to_signed(1, 8),
    to_signed(2, 8),
    to_signed(4, 8),
    to_signed(5, 8),
    to_signed(5, 8),
    to_signed(3, 8),
    to_signed(0, 8),
    to_signed(-4, 8),
    to_signed(-7, 8),
    to_signed(-10, 8),
    to_signed(-10, 8),
    to_signed(-7, 8),
    to_signed(-3, 8),
    to_signed(0, 8),
    to_signed(2, 8),
    to_signed(2, 8),
    to_signed(2, 8),
    to_signed(2, 8),
    to_signed(3, 8),
    to_signed(3, 8),
    to_signed(3, 8),
    to_signed(2, 8),
    to_signed(4, 8),
    to_signed(7, 8),
    to_signed(9, 8),
    to_signed(10, 8),
    to_signed(10, 8),
    to_signed(8, 8),
    to_signed(6, 8),
    to_signed(4, 8),
    to_signed(3, 8),
    to_signed(3, 8),
    to_signed(3, 8),
    to_signed(4, 8),
    to_signed(5, 8),
    to_signed(6, 8),
    to_signed(7, 8),
    to_signed(8, 8),
    to_signed(9, 8),
    to_signed(9, 8),
    to_signed(9, 8),
    to_signed(7, 8),
    to_signed(5, 8),
    to_signed(4, 8),
    to_signed(3, 8),
    to_signed(3, 8),
    to_signed(3, 8),
    to_signed(4, 8),
    to_signed(3, 8),
    to_signed(1, 8),
    to_signed(-1, 8),
    to_signed(-2, 8),
    to_signed(-4, 8),
    to_signed(-4, 8),
    to_signed(-4, 8),
    to_signed(-3, 8),
    to_signed(-2, 8),
    to_signed(-1, 8),
    to_signed(-1, 8),
    to_signed(0, 8),
    to_signed(1, 8),
    to_signed(0, 8),
    to_signed(-2, 8),
    to_signed(-4, 8),
    to_signed(-5, 8),
    to_signed(-5, 8),
    to_signed(-4, 8),
    to_signed(-2, 8),
    to_signed(1, 8),
    to_signed(3, 8),
    to_signed(3, 8),
    to_signed(2, 8),
    to_signed(1, 8),
    to_signed(1, 8),
    to_signed(-1, 8),
    to_signed(-2, 8),
    to_signed(-2, 8),
    to_signed(-1, 8),
    to_signed(0, 8),
    to_signed(1, 8),
    to_signed(3, 8),
    to_signed(7, 8),
    to_signed(9, 8),
    to_signed(9, 8),
    to_signed(6, 8),
    to_signed(4, 8),
    to_signed(3, 8),
    to_signed(2, 8),
    to_signed(3, 8),
    to_signed(5, 8),
    to_signed(7, 8),
    to_signed(8, 8),
    to_signed(7, 8),
    to_signed(6, 8),
    to_signed(5, 8),
    to_signed(4, 8),
    to_signed(2, 8),
    to_signed(-1, 8),
    to_signed(-3, 8),
    to_signed(-4, 8),
    to_signed(-4, 8),
    to_signed(-4, 8),
    to_signed(-3, 8),
    to_signed(-2, 8),
    to_signed(0, 8),
    to_signed(1, 8),
    to_signed(1, 8),
    to_signed(0, 8),
    to_signed(-1, 8),
    to_signed(-2, 8),
    to_signed(-5, 8),
    to_signed(-7, 8),
    to_signed(-8, 8),
    to_signed(-7, 8),
    to_signed(-6, 8),
    to_signed(-5, 8),
    to_signed(-4, 8),
    to_signed(-4, 8),
    to_signed(-5, 8),
    to_signed(-7, 8),
    to_signed(-10, 8),
    to_signed(-12, 8),
    to_signed(-13, 8),
    to_signed(-13, 8),
    to_signed(-12, 8),
    to_signed(-10, 8),
    to_signed(-7, 8),
    to_signed(-5, 8),
    to_signed(-4, 8),
    to_signed(-3, 8),
    to_signed(-2, 8),
    to_signed(-2, 8),
    to_signed(-2, 8),
    to_signed(-1, 8),
    to_signed(0, 8),
    to_signed(0, 8),
    to_signed(1, 8),
    to_signed(1, 8),
    to_signed(2, 8),
    to_signed(1, 8),
    to_signed(0, 8),
    to_signed(-1, 8),
    to_signed(-3, 8),
    to_signed(-5, 8),
    to_signed(-6, 8),
    to_signed(-6, 8),
    to_signed(-4, 8),
    to_signed(-1, 8),
    to_signed(1, 8),
    to_signed(3, 8),
    to_signed(6, 8),
    to_signed(7, 8),
    to_signed(7, 8),
    to_signed(7, 8),
    to_signed(6, 8),
    to_signed(5, 8),
    to_signed(3, 8),
    to_signed(3, 8),
    to_signed(5, 8),
    to_signed(6, 8),
    to_signed(6, 8),
    to_signed(3, 8),
    to_signed(1, 8),
    to_signed(-2, 8),
    to_signed(-5, 8),
    to_signed(-8, 8),
    to_signed(-11, 8),
    to_signed(-12, 8),
    to_signed(-10, 8),
    to_signed(-6, 8),
    to_signed(-3, 8),
    to_signed(-1, 8),
    to_signed(-1, 8),
    to_signed(-2, 8),
    to_signed(-3, 8),
    to_signed(-5, 8),
    to_signed(-6, 8),
    to_signed(-6, 8),
    to_signed(-7, 8),
    to_signed(-8, 8),
    to_signed(-9, 8),
    to_signed(-8, 8),
    to_signed(-7, 8),
    to_signed(-7, 8),
    to_signed(-6, 8),
    to_signed(-7, 8),
    to_signed(-8, 8),
    to_signed(-11, 8),
    to_signed(-13, 8),
    to_signed(-13, 8),
    to_signed(-11, 8),
    to_signed(-8, 8),
    to_signed(-5, 8),
    to_signed(-3, 8),
    to_signed(-1, 8),
    to_signed(2, 8),
    to_signed(4, 8),
    to_signed(4, 8),
    to_signed(3, 8),
    to_signed(2, 8),
    to_signed(1, 8),
    to_signed(0, 8),
    to_signed(-1, 8),
    to_signed(-1, 8),
    to_signed(-1, 8),
    to_signed(1, 8),
    to_signed(3, 8),
    to_signed(4, 8),
    to_signed(3, 8),
    to_signed(1, 8),
    to_signed(-1, 8),
    to_signed(-2, 8),
    to_signed(-3, 8),
    to_signed(-2, 8),
    to_signed(1, 8),
    to_signed(4, 8),
    to_signed(4, 8),
    to_signed(3, 8),
    to_signed(2, 8),
    to_signed(1, 8),
    to_signed(0, 8),
    to_signed(-1, 8),
    to_signed(-2, 8),
    to_signed(-4, 8),
    to_signed(-5, 8),
    to_signed(-6, 8),
    to_signed(-6, 8),
    to_signed(-5, 8),
    to_signed(-4, 8),
    to_signed(-3, 8),
    to_signed(-4, 8),
    to_signed(-7, 8),
    to_signed(-10, 8),
    to_signed(-11, 8),
    to_signed(-10, 8),
    to_signed(-6, 8),
    to_signed(-3, 8),
    to_signed(-1, 8),
    to_signed(-1, 8),
    to_signed(-1, 8),
    to_signed(-2, 8),
    to_signed(-4, 8),
    to_signed(-5, 8),
    to_signed(-5, 8),
    to_signed(-5, 8),
    to_signed(-5, 8),
    to_signed(-6, 8),
    to_signed(-7, 8),
    to_signed(-8, 8),
    to_signed(-9, 8),
    to_signed(-8, 8),
    to_signed(-7, 8),
    to_signed(-6, 8),
    to_signed(-6, 8),
    to_signed(-6, 8),
    to_signed(-5, 8),
    to_signed(-4, 8),
    to_signed(-1, 8),
    to_signed(2, 8),
    to_signed(4, 8),
    to_signed(6, 8),
    to_signed(7, 8),
    to_signed(8, 8),
    to_signed(9, 8),
    to_signed(10, 8),
    to_signed(11, 8),
    to_signed(12, 8),
    to_signed(12, 8),
    to_signed(11, 8),
    to_signed(9, 8),
    to_signed(8, 8),
    to_signed(9, 8),
    to_signed(10, 8),
    to_signed(9, 8),
    to_signed(7, 8),
    to_signed(5, 8),
    to_signed(3, 8),
    to_signed(1, 8),
    to_signed(0, 8),
    to_signed(0, 8),
    to_signed(2, 8),
    to_signed(4, 8),
    to_signed(5, 8),
    to_signed(6, 8),
    to_signed(5, 8),
    to_signed(4, 8),
    to_signed(4, 8),
    to_signed(5, 8),
    to_signed(6, 8),
    to_signed(7, 8),
    to_signed(6, 8),
    to_signed(5, 8),
    to_signed(3, 8),
    to_signed(1, 8),
    to_signed(-3, 8),
    to_signed(-7, 8),
    to_signed(-10, 8),
    to_signed(-12, 8),
    to_signed(-12, 8),
    to_signed(-11, 8),
    to_signed(-11, 8),
    to_signed(-10, 8),
    to_signed(-8, 8),
    to_signed(-5, 8),
    to_signed(-3, 8),
    to_signed(-1, 8),
    to_signed(1, 8),
    to_signed(2, 8),
    to_signed(3, 8),
    to_signed(5, 8),
    to_signed(6, 8),
    to_signed(7, 8),
    to_signed(8, 8),
    to_signed(7, 8),
    to_signed(5, 8),
    to_signed(3, 8),
    to_signed(2, 8),
    to_signed(1, 8),
    to_signed(0, 8),
    to_signed(-1, 8),
    to_signed(-3, 8),
    to_signed(-4, 8),
    to_signed(-4, 8),
    to_signed(-2, 8),
    to_signed(-1, 8),
    to_signed(1, 8),
    to_signed(2, 8),
    to_signed(2, 8),
    to_signed(1, 8),
    to_signed(0, 8),
    to_signed(-1, 8),
    to_signed(1, 8),
    to_signed(2, 8),
    to_signed(3, 8),
    to_signed(2, 8),
    to_signed(1, 8),
    to_signed(0, 8),
    to_signed(-1, 8),
    to_signed(-3, 8),
    to_signed(-4, 8),
    to_signed(-4, 8),
    to_signed(-4, 8),
    to_signed(-4, 8),
    to_signed(-3, 8),
    to_signed(-2, 8),
    to_signed(-1, 8),
    to_signed(0, 8),
    to_signed(1, 8),
    to_signed(2, 8),
    to_signed(2, 8),
    to_signed(1, 8),
    to_signed(0, 8),
    to_signed(-1, 8),
    to_signed(0, 8),
    to_signed(1, 8),
    to_signed(3, 8),
    to_signed(2, 8),
    to_signed(1, 8),
    to_signed(1, 8),
    to_signed(1, 8),
    to_signed(0, 8),
    to_signed(-3, 8),
    to_signed(-4, 8),
    to_signed(-4, 8),
    to_signed(-2, 8),
    to_signed(0, 8),
    to_signed(2, 8),
    to_signed(3, 8),
    to_signed(6, 8),
    to_signed(8, 8),
    to_signed(8, 8),
    to_signed(6, 8),
    to_signed(3, 8),
    to_signed(1, 8),
    to_signed(1, 8),
    to_signed(2, 8),
    to_signed(3, 8),
    to_signed(4, 8),
    to_signed(4, 8),
    to_signed(3, 8),
    to_signed(1, 8),
    to_signed(-2, 8),
    to_signed(-4, 8),
    to_signed(-6, 8),
    to_signed(-6, 8),
    to_signed(-4, 8),
    to_signed(-2, 8),
    to_signed(-1, 8),
    to_signed(0, 8),
    to_signed(1, 8),
    to_signed(1, 8),
    to_signed(1, 8),
    to_signed(-1, 8),
    to_signed(-3, 8),
    to_signed(-5, 8),
    to_signed(-5, 8),
    to_signed(-5, 8),
    to_signed(-4, 8),
    to_signed(-4, 8),
    to_signed(-3, 8),
    to_signed(-4, 8),
    to_signed(-5, 8),
    to_signed(-7, 8),
    to_signed(-9, 8),
    to_signed(-10, 8),
    to_signed(-11, 8),
    to_signed(-12, 8),
    to_signed(-13, 8),
    to_signed(-12, 8),
    to_signed(-10, 8),
    to_signed(-8, 8),
    to_signed(-5, 8),
    to_signed(-2, 8),
    to_signed(-1, 8),
    to_signed(-1, 8),
    to_signed(-2, 8),
    to_signed(-2, 8),
    to_signed(-2, 8),
    to_signed(-1, 8),
    to_signed(1, 8),
    to_signed(4, 8),
    to_signed(6, 8),
    to_signed(6, 8),
    to_signed(5, 8),
    to_signed(3, 8),
    to_signed(1, 8),
    to_signed(-1, 8),
    to_signed(-2, 8),
    to_signed(-3, 8),
    to_signed(-4, 8),
    to_signed(-4, 8),
    to_signed(-3, 8),
    to_signed(-1, 8),
    to_signed(1, 8),
    to_signed(4, 8),
    to_signed(6, 8),
    to_signed(6, 8),
    to_signed(5, 8),
    to_signed(4, 8),
    to_signed(4, 8),
    to_signed(6, 8),
    to_signed(10, 8),
    to_signed(13, 8),
    to_signed(15, 8),
    to_signed(14, 8),
    to_signed(13, 8),
    to_signed(12, 8),
    to_signed(9, 8),
    to_signed(5, 8),
    to_signed(0, 8),
    to_signed(-3, 8),
    to_signed(-5, 8),
    to_signed(-5, 8),
    to_signed(-4, 8),
    to_signed(-3, 8),
    to_signed(-1, 8),
    to_signed(0, 8),
    to_signed(0, 8),
    to_signed(0, 8),
    to_signed(-2, 8),
    to_signed(-3, 8),
    to_signed(-3, 8),
    to_signed(-1, 8),
    to_signed(1, 8),
    to_signed(4, 8),
    to_signed(6, 8),
    to_signed(6, 8),
    to_signed(4, 8),
    to_signed(1, 8),
    to_signed(-2, 8),
    to_signed(-5, 8),
    to_signed(-8, 8),
    to_signed(-10, 8),
    to_signed(-11, 8),
    to_signed(-11, 8),
    to_signed(-10, 8),
    to_signed(-9, 8),
    to_signed(-6, 8),
    to_signed(-4, 8),
    to_signed(-3, 8),
    to_signed(-2, 8),
    to_signed(-2, 8),
    to_signed(-1, 8),
    to_signed(-1, 8),
    to_signed(-1, 8),
    to_signed(-1, 8),
    to_signed(1, 8),
    to_signed(4, 8),
    to_signed(5, 8),
    to_signed(5, 8),
    to_signed(4, 8),
    to_signed(4, 8),
    to_signed(3, 8),
    to_signed(1, 8),
    to_signed(-1, 8),
    to_signed(-2, 8),
    to_signed(-2, 8),
    to_signed(2, 8),
    to_signed(6, 8),
    to_signed(9, 8),
    to_signed(11, 8),
    to_signed(11, 8),
    to_signed(9, 8),
    to_signed(7, 8),
    to_signed(4, 8),
    to_signed(3, 8),
    to_signed(3, 8),
    to_signed(3, 8),
    to_signed(3, 8),
    to_signed(3, 8),
    to_signed(3, 8),
    to_signed(2, 8),
    to_signed(1, 8),
    to_signed(0, 8),
    to_signed(-1, 8),
    to_signed(-3, 8),
    to_signed(-7, 8),
    to_signed(-9, 8),
    to_signed(-9, 8),
    to_signed(-6, 8),
    to_signed(-4, 8),
    to_signed(-3, 8),
    to_signed(-3, 8),
    to_signed(-2, 8),
    to_signed(-3, 8),
    to_signed(-4, 8),
    to_signed(-6, 8),
    to_signed(-7, 8),
    to_signed(-7, 8),
    to_signed(-7, 8),
    to_signed(-7, 8),
    to_signed(-7, 8),
    to_signed(-6, 8),
    to_signed(-6, 8),
    to_signed(-6, 8),
    to_signed(-6, 8),
    to_signed(-7, 8),
    to_signed(-7, 8),
    to_signed(-8, 8),
    to_signed(-9, 8),
    to_signed(-8, 8),
    to_signed(-5, 8),
    to_signed(-1, 8),
    to_signed(3, 8),
    to_signed(6, 8),
    to_signed(8, 8),
    to_signed(8, 8),
    to_signed(5, 8),
    to_signed(2, 8),
    to_signed(0, 8),
    to_signed(-1, 8),
    to_signed(1, 8),
    to_signed(4, 8),
    to_signed(6, 8),
    to_signed(6, 8),
    to_signed(5, 8),
    to_signed(3, 8),
    to_signed(1, 8),
    to_signed(-2, 8),
    to_signed(-4, 8),
    to_signed(-7, 8),
    to_signed(-9, 8),
    to_signed(-9, 8),
    to_signed(-7, 8),
    to_signed(-4, 8),
    to_signed(-1, 8),
    to_signed(2, 8),
    to_signed(4, 8),
    to_signed(4, 8),
    to_signed(2, 8),
    to_signed(0, 8),
    to_signed(-1, 8),
    to_signed(-2, 8),
    to_signed(-1, 8),
    to_signed(3, 8),
    to_signed(7, 8),
    to_signed(8, 8),
    to_signed(7, 8),
    to_signed(4, 8),
    to_signed(1, 8),
    to_signed(-2, 8),
    to_signed(-5, 8),
    to_signed(-9, 8),
    to_signed(-12, 8),
    to_signed(-14, 8),
    to_signed(-13, 8),
    to_signed(-9, 8),
    to_signed(-7, 8),
    to_signed(-5, 8),
    to_signed(-4, 8),
    to_signed(-4, 8),
    to_signed(-5, 8),
    to_signed(-6, 8),
    to_signed(-7, 8),
    to_signed(-7, 8),
    to_signed(-6, 8),
    to_signed(-3, 8),
    to_signed(0, 8),
    to_signed(3, 8),
    to_signed(4, 8),
    to_signed(4, 8),
    to_signed(1, 8),
    to_signed(-3, 8),
    to_signed(-8, 8),
    to_signed(-12, 8),
    to_signed(-13, 8),
    to_signed(-11, 8),
    to_signed(-9, 8),
    to_signed(-6, 8),
    to_signed(-3, 8),
    to_signed(0, 8),
    to_signed(2, 8),
    to_signed(3, 8),
    to_signed(2, 8),
    to_signed(1, 8),
    to_signed(-1, 8),
    to_signed(-1, 8),
    to_signed(2, 8),
    to_signed(6, 8),
    to_signed(10, 8),
    to_signed(12, 8),
    to_signed(13, 8),
    to_signed(13, 8),
    to_signed(10, 8),
    to_signed(6, 8),
    to_signed(2, 8),
    to_signed(-1, 8),
    to_signed(-3, 8),
    to_signed(-3, 8),
    to_signed(0, 8),
    to_signed(4, 8),
    to_signed(7, 8),
    to_signed(9, 8),
    to_signed(9, 8),
    to_signed(7, 8),
    to_signed(5, 8),
    to_signed(3, 8),
    to_signed(2, 8),
    to_signed(1, 8),
    to_signed(3, 8),
    to_signed(4, 8),
    to_signed(4, 8),
    to_signed(5, 8),
    to_signed(6, 8),
    to_signed(7, 8),
    to_signed(6, 8),
    to_signed(4, 8),
    to_signed(-1, 8),
    to_signed(-5, 8),
    to_signed(-8, 8),
    to_signed(-7, 8),
    to_signed(-4, 8),
    to_signed(0, 8),
    to_signed(3, 8),
    to_signed(5, 8),
    to_signed(6, 8),
    to_signed(5, 8),
    to_signed(4, 8),
    to_signed(1, 8),
    to_signed(-1, 8),
    to_signed(-4, 8),
    to_signed(-6, 8),
    to_signed(-5, 8),
    to_signed(-2, 8),
    to_signed(0, 8),
    to_signed(1, 8),
    to_signed(1, 8),
    to_signed(0, 8),
    to_signed(-1, 8),
    to_signed(-4, 8),
    to_signed(-7, 8),
    to_signed(-8, 8),
    to_signed(-8, 8),
    to_signed(-4, 8),
    to_signed(0, 8),
    to_signed(5, 8),
    to_signed(8, 8),
    to_signed(10, 8),
    to_signed(10, 8),
    to_signed(8, 8),
    to_signed(6, 8),
    to_signed(3, 8),
    to_signed(2, 8),
    to_signed(3, 8),
    to_signed(5, 8),
    to_signed(7, 8),
    to_signed(8, 8),
    to_signed(8, 8),
    to_signed(7, 8),
    to_signed(7, 8),
    to_signed(7, 8),
    to_signed(6, 8),
    to_signed(4, 8),
    to_signed(1, 8),
    to_signed(0, 8),
    to_signed(1, 8),
    to_signed(4, 8),
    to_signed(8, 8),
    to_signed(11, 8),
    to_signed(13, 8),
    to_signed(13, 8),
    to_signed(12, 8),
    to_signed(9, 8),
    to_signed(6, 8),
    to_signed(4, 8),
    to_signed(4, 8),
    to_signed(5, 8),
    to_signed(7, 8),
    to_signed(10, 8),
    to_signed(11, 8),
    to_signed(9, 8),
    to_signed(6, 8),
    to_signed(4, 8),
    to_signed(2, 8),
    to_signed(0, 8),
    to_signed(-1, 8),
    to_signed(-2, 8),
    to_signed(-1, 8),
    to_signed(1, 8),
    to_signed(4, 8),
    to_signed(7, 8),
    to_signed(8, 8),
    to_signed(8, 8),
    to_signed(7, 8),
    to_signed(6, 8),
    to_signed(4, 8),
    to_signed(3, 8),
    to_signed(4, 8),
    to_signed(7, 8),
    to_signed(9, 8),
    to_signed(10, 8),
    to_signed(8, 8),
    to_signed(6, 8),
    to_signed(3, 8),
    to_signed(0, 8),
    to_signed(-2, 8),
    to_signed(-3, 8),
    to_signed(-5, 8),
    to_signed(-7, 8),
    to_signed(-7, 8),
    to_signed(-6, 8),
    to_signed(-4, 8),
    to_signed(-3, 8),
    to_signed(-2, 8),
    to_signed(-2, 8),
    to_signed(-2, 8),
    to_signed(-1, 8),
    to_signed(-1, 8),
    to_signed(-1, 8),
    to_signed(0, 8),
    to_signed(2, 8),
    to_signed(4, 8),
    to_signed(4, 8),
    to_signed(3, 8),
    to_signed(2, 8),
    to_signed(0, 8),
    to_signed(-3, 8),
    to_signed(-6, 8),
    to_signed(-9, 8),
    to_signed(-10, 8),
    to_signed(-10, 8),
    to_signed(-8, 8),
    to_signed(-5, 8),
    to_signed(-2, 8),
    to_signed(0, 8),
    to_signed(1, 8),
    to_signed(2, 8),
    to_signed(1, 8),
    to_signed(1, 8),
    to_signed(1, 8),
    to_signed(2, 8),
    to_signed(2, 8),
    to_signed(3, 8),
    to_signed(5, 8),
    to_signed(7, 8),
    to_signed(7, 8),
    to_signed(6, 8),
    to_signed(4, 8),
    to_signed(1, 8),
    to_signed(-3, 8),
    to_signed(-6, 8),
    to_signed(-9, 8),
    to_signed(-9, 8),
    to_signed(-7, 8),
    to_signed(-4, 8),
    to_signed(-1, 8),
    to_signed(1, 8),
    to_signed(2, 8),
    to_signed(0, 8),
    to_signed(-3, 8),
    to_signed(-5, 8),
    to_signed(-6, 8),
    to_signed(-6, 8),
    to_signed(-6, 8),
    to_signed(-5, 8),
    to_signed(-5, 8),
    to_signed(-4, 8),
    to_signed(-4, 8),
    to_signed(-5, 8),
    to_signed(-7, 8),
    to_signed(-9, 8),
    to_signed(-10, 8),
    to_signed(-12, 8),
    to_signed(-14, 8),
    to_signed(-15, 8),
    to_signed(-13, 8),
    to_signed(-7, 8),
    to_signed(-2, 8),
    to_signed(0, 8),
    to_signed(0, 8),
    to_signed(-1, 8),
    to_signed(-2, 8),
    to_signed(-4, 8),
    to_signed(-5, 8),
    to_signed(-6, 8),
    to_signed(-5, 8),
    to_signed(-4, 8),
    to_signed(-2, 8),
    to_signed(-1, 8),
    to_signed(1, 8),
    to_signed(2, 8),
    to_signed(1, 8),
    to_signed(-1, 8),
    to_signed(-3, 8),
    to_signed(-6, 8),
    to_signed(-7, 8),
    to_signed(-7, 8),
    to_signed(-5, 8),
    to_signed(0, 8),
    to_signed(5, 8),
    to_signed(9, 8),
    to_signed(11, 8),
    to_signed(11, 8),
    to_signed(8, 8),
    to_signed(5, 8),
    to_signed(2, 8),
    to_signed(0, 8),
    to_signed(0, 8),
    to_signed(2, 8),
    to_signed(4, 8),
    to_signed(6, 8),
    to_signed(6, 8),
    to_signed(5, 8),
    to_signed(2, 8),
    to_signed(-2, 8),
    to_signed(-5, 8),
    to_signed(-7, 8),
    to_signed(-8, 8),
    to_signed(-8, 8),
    to_signed(-5, 8),
    to_signed(-3, 8),
    to_signed(0, 8),
    to_signed(0, 8),
    to_signed(-2, 8),
    to_signed(-4, 8),
    to_signed(-7, 8),
    to_signed(-10, 8),
    to_signed(-11, 8),
    to_signed(-12, 8),
    to_signed(-11, 8),
    to_signed(-8, 8),
    to_signed(-6, 8),
    to_signed(-4, 8),
    to_signed(-4, 8),
    to_signed(-6, 8),
    to_signed(-9, 8),
    to_signed(-13, 8),
    to_signed(-18, 8),
    to_signed(-20, 8),
    to_signed(-20, 8),
    to_signed(-18, 8),
    to_signed(-15, 8),
    to_signed(-11, 8),
    to_signed(-7, 8),
    to_signed(-4, 8),
    to_signed(-3, 8),
    to_signed(-3, 8),
    to_signed(-4, 8),
    to_signed(-5, 8),
    to_signed(-6, 8),
    to_signed(-5, 8),
    to_signed(-2, 8),
    to_signed(2, 8),
    to_signed(6, 8),
    to_signed(9, 8),
    to_signed(11, 8),
    to_signed(9, 8),
    to_signed(7, 8),
    to_signed(5, 8),
    to_signed(3, 8),
    to_signed(1, 8),
    to_signed(0, 8),
    to_signed(1, 8),
    to_signed(2, 8),
    to_signed(3, 8),
    to_signed(5, 8),
    to_signed(7, 8),
    to_signed(8, 8),
    to_signed(7, 8),
    to_signed(6, 8),
    to_signed(4, 8),
    to_signed(3, 8),
    to_signed(3, 8),
    to_signed(3, 8),
    to_signed(4, 8),
    to_signed(4, 8),
    to_signed(5, 8),
    to_signed(5, 8),
    to_signed(3, 8),
    to_signed(-1, 8),
    to_signed(-3, 8),
    to_signed(-6, 8),
    to_signed(-9, 8),
    to_signed(-11, 8),
    to_signed(-11, 8),
    to_signed(-9, 8),
    to_signed(-7, 8),
    to_signed(-5, 8),
    to_signed(-5, 8),
    to_signed(-7, 8),
    to_signed(-10, 8),
    to_signed(-12, 8),
    to_signed(-11, 8),
    to_signed(-9, 8),
    to_signed(-6, 8),
    to_signed(-3, 8),
    to_signed(-1, 8),
    to_signed(0, 8),
    to_signed(0, 8),
    to_signed(-2, 8),
    to_signed(-5, 8),
    to_signed(-8, 8),
    to_signed(-12, 8),
    to_signed(-13, 8),
    to_signed(-14, 8),
    to_signed(-13, 8),
    to_signed(-11, 8),
    to_signed(-7, 8),
    to_signed(-4, 8),
    to_signed(-2, 8),
    to_signed(-2, 8),
    to_signed(-2, 8),
    to_signed(-5, 8),
    to_signed(-8, 8),
    to_signed(-10, 8),
    to_signed(-9, 8),
    to_signed(-6, 8),
    to_signed(-2, 8),
    to_signed(3, 8),
    to_signed(7, 8),
    to_signed(9, 8),
    to_signed(9, 8),
    to_signed(6, 8),
    to_signed(2, 8),
    to_signed(-2, 8),
    to_signed(-6, 8),
    to_signed(-8, 8),
    to_signed(-7, 8),
    to_signed(-3, 8),
    to_signed(3, 8),
    to_signed(8, 8),
    to_signed(12, 8),
    to_signed(13, 8),
    to_signed(10, 8),
    to_signed(5, 8),
    to_signed(0, 8),
    to_signed(-3, 8),
    to_signed(-4, 8),
    to_signed(-4, 8),
    to_signed(-3, 8),
    to_signed(-1, 8),
    to_signed(2, 8),
    to_signed(3, 8),
    to_signed(3, 8),
    to_signed(0, 8),
    to_signed(-3, 8),
    to_signed(-7, 8),
    to_signed(-11, 8),
    to_signed(-15, 8),
    to_signed(-15, 8),
    to_signed(-12, 8),
    to_signed(-8, 8),
    to_signed(-5, 8),
    to_signed(-2, 8),
    to_signed(0, 8),
    to_signed(0, 8),
    to_signed(-1, 8),
    to_signed(-4, 8),
    to_signed(-7, 8),
    to_signed(-9, 8),
    to_signed(-8, 8),
    to_signed(-4, 8),
    to_signed(0, 8),
    to_signed(4, 8),
    to_signed(6, 8),
    to_signed(5, 8),
    to_signed(2, 8),
    to_signed(-2, 8),
    to_signed(-5, 8),
    to_signed(-6, 8),
    to_signed(-6, 8),
    to_signed(-4, 8),
    to_signed(-1, 8),
    to_signed(3, 8),
    to_signed(6, 8),
    to_signed(8, 8),
    to_signed(9, 8),
    to_signed(8, 8),
    to_signed(5, 8),
    to_signed(3, 8),
    to_signed(3, 8),
    to_signed(4, 8),
    to_signed(6, 8),
    to_signed(9, 8),
    to_signed(12, 8),
    to_signed(14, 8),
    to_signed(12, 8),
    to_signed(9, 8),
    to_signed(4, 8),
    to_signed(1, 8),
    to_signed(-3, 8),
    to_signed(-6, 8),
    to_signed(-8, 8),
    to_signed(-8, 8),
    to_signed(-5, 8),
    to_signed(-2, 8),
    to_signed(0, 8),
    to_signed(1, 8),
    to_signed(2, 8),
    to_signed(1, 8),
    to_signed(-2, 8),
    to_signed(-5, 8),
    to_signed(-6, 8),
    to_signed(-5, 8),
    to_signed(-2, 8),
    to_signed(1, 8),
    to_signed(6, 8),
    to_signed(10, 8),
    to_signed(11, 8),
    to_signed(9, 8),
    to_signed(3, 8),
    to_signed(-3, 8),
    to_signed(-8, 8),
    to_signed(-12, 8),
    to_signed(-14, 8),
    to_signed(-15, 8),
    to_signed(-13, 8),
    to_signed(-12, 8),
    to_signed(-9, 8),
    to_signed(-6, 8),
    to_signed(-4, 8),
    to_signed(-5, 8),
    to_signed(-8, 8),
    to_signed(-10, 8),
    to_signed(-11, 8),
    to_signed(-11, 8),
    to_signed(-8, 8),
    to_signed(-3, 8),
    to_signed(3, 8),
    to_signed(7, 8),
    to_signed(9, 8),
    to_signed(8, 8),
    to_signed(5, 8),
    to_signed(1, 8),
    to_signed(-4, 8),
    to_signed(-7, 8),
    to_signed(-7, 8),
    to_signed(-5, 8),
    to_signed(-2, 8),
    to_signed(3, 8),
    to_signed(7, 8),
    to_signed(9, 8),
    to_signed(9, 8),
    to_signed(8, 8),
    to_signed(5, 8),
    to_signed(3, 8),
    to_signed(2, 8),
    to_signed(2, 8),
    to_signed(6, 8),
    to_signed(11, 8),
    to_signed(16, 8),
    to_signed(20, 8),
    to_signed(20, 8),
    to_signed(18, 8),
    to_signed(13, 8),
    to_signed(7, 8),
    to_signed(1, 8),
    to_signed(-3, 8),
    to_signed(-4, 8),
    to_signed(-2, 8),
    to_signed(2, 8),
    to_signed(6, 8),
    to_signed(9, 8),
    to_signed(10, 8),
    to_signed(10, 8),
    to_signed(6, 8),
    to_signed(-1, 8),
    to_signed(-7, 8),
    to_signed(-10, 8),
    to_signed(-10, 8),
    to_signed(-8, 8),
    to_signed(-3, 8),
    to_signed(2, 8),
    to_signed(6, 8),
    to_signed(7, 8),
    to_signed(5, 8),
    to_signed(1, 8),
    to_signed(-4, 8),
    to_signed(-10, 8),
    to_signed(-13, 8),
    to_signed(-13, 8),
    to_signed(-10, 8),
    to_signed(-5, 8),
    to_signed(1, 8),
    to_signed(5, 8),
    to_signed(8, 8),
    to_signed(6, 8),
    to_signed(2, 8),
    to_signed(-2, 8),
    to_signed(-6, 8),
    to_signed(-9, 8),
    to_signed(-9, 8),
    to_signed(-6, 8),
    to_signed(0, 8),
    to_signed(4, 8),
    to_signed(5, 8),
    to_signed(6, 8),
    to_signed(5, 8),
    to_signed(2, 8),
    to_signed(-2, 8),
    to_signed(-6, 8),
    to_signed(-8, 8),
    to_signed(-8, 8),
    to_signed(-6, 8),
    to_signed(0, 8),
    to_signed(5, 8),
    to_signed(10, 8),
    to_signed(13, 8),
    to_signed(13, 8),
    to_signed(10, 8),
    to_signed(6, 8),
    to_signed(2, 8),
    to_signed(0, 8),
    to_signed(-1, 8),
    to_signed(2, 8),
    to_signed(7, 8),
    to_signed(11, 8),
    to_signed(13, 8),
    to_signed(13, 8),
    to_signed(10, 8),
    to_signed(6, 8),
    to_signed(1, 8),
    to_signed(-2, 8),
    to_signed(-4, 8),
    to_signed(-4, 8),
    to_signed(-3, 8),
    to_signed(0, 8),
    to_signed(2, 8),
    to_signed(4, 8),
    to_signed(5, 8),
    to_signed(3, 8),
    to_signed(-1, 8),
    to_signed(-6, 8),
    to_signed(-8, 8),
    to_signed(-9, 8),
    to_signed(-9, 8),
    to_signed(-6, 8),
    to_signed(-1, 8),
    to_signed(3, 8),
    to_signed(3, 8),
    to_signed(1, 8),
    to_signed(-2, 8),
    to_signed(-6, 8),
    to_signed(-12, 8),
    to_signed(-16, 8),
    to_signed(-18, 8),
    to_signed(-17, 8),
    to_signed(-16, 8),
    to_signed(-14, 8),
    to_signed(-10, 8),
    to_signed(-7, 8),
    to_signed(-6, 8),
    to_signed(-6, 8),
    to_signed(-8, 8),
    to_signed(-9, 8),
    to_signed(-10, 8),
    to_signed(-10, 8),
    to_signed(-9, 8),
    to_signed(-6, 8),
    to_signed(-1, 8),
    to_signed(4, 8),
    to_signed(8, 8),
    to_signed(8, 8),
    to_signed(7, 8),
    to_signed(4, 8),
    to_signed(1, 8),
    to_signed(-2, 8),
    to_signed(-3, 8),
    to_signed(-3, 8),
    to_signed(-2, 8),
    to_signed(0, 8),
    to_signed(1, 8),
    to_signed(3, 8),
    to_signed(5, 8),
    to_signed(5, 8),
    to_signed(4, 8),
    to_signed(2, 8),
    to_signed(2, 8),
    to_signed(1, 8),
    to_signed(1, 8),
    to_signed(4, 8),
    to_signed(8, 8),
    to_signed(11, 8),
    to_signed(13, 8),
    to_signed(14, 8),
    to_signed(11, 8),
    to_signed(7, 8),
    to_signed(1, 8),
    to_signed(-2, 8),
    to_signed(-4, 8),
    to_signed(-4, 8),
    to_signed(-2, 8),
    to_signed(2, 8),
    to_signed(5, 8),
    to_signed(6, 8),
    to_signed(6, 8),
    to_signed(4, 8),
    to_signed(0, 8),
    to_signed(-2, 8),
    to_signed(-3, 8),
    to_signed(-2, 8),
    to_signed(1, 8),
    to_signed(3, 8),
    to_signed(5, 8),
    to_signed(6, 8),
    to_signed(7, 8),
    to_signed(6, 8),
    to_signed(3, 8),
    to_signed(-3, 8),
    to_signed(-7, 8),
    to_signed(-10, 8),
    to_signed(-12, 8),
    to_signed(-12, 8),
    to_signed(-10, 8),
    to_signed(-6, 8),
    to_signed(-2, 8),
    to_signed(0, 8),
    to_signed(0, 8),
    to_signed(-1, 8),
    to_signed(-4, 8),
    to_signed(-7, 8),
    to_signed(-10, 8),
    to_signed(-12, 8),
    to_signed(-12, 8),
    to_signed(-10, 8),
    to_signed(-6, 8),
    to_signed(-1, 8),
    to_signed(2, 8),
    to_signed(4, 8),
    to_signed(5, 8),
    to_signed(4, 8),
    to_signed(1, 8),
    to_signed(-3, 8),
    to_signed(-6, 8),
    to_signed(-7, 8),
    to_signed(-6, 8),
    to_signed(-2, 8),
    to_signed(3, 8),
    to_signed(9, 8),
    to_signed(13, 8),
    to_signed(13, 8),
    to_signed(10, 8),
    to_signed(7, 8),
    to_signed(4, 8),
    to_signed(2, 8),
    to_signed(2, 8),
    to_signed(2, 8),
    to_signed(2, 8),
    to_signed(1, 8),
    to_signed(4, 8),
    to_signed(8, 8),
    to_signed(9, 8),
    to_signed(8, 8),
    to_signed(6, 8),
    to_signed(3, 8),
    to_signed(-2, 8),
    to_signed(-6, 8),
    to_signed(-7, 8),
    to_signed(-5, 8),
    to_signed(-3, 8),
    to_signed(-1, 8),
    to_signed(1, 8),
    to_signed(2, 8),
    to_signed(1, 8),
    to_signed(-2, 8),
    to_signed(-3, 8),
    to_signed(-3, 8),
    to_signed(-3, 8),
    to_signed(-2, 8),
    to_signed(-1, 8),
    to_signed(1, 8),
    to_signed(2, 8),
    to_signed(2, 8),
    to_signed(3, 8),
    to_signed(3, 8),
    to_signed(3, 8),
    to_signed(1, 8),
    to_signed(-1, 8),
    to_signed(-3, 8),
    to_signed(-3, 8),
    to_signed(-2, 8),
    to_signed(0, 8),
    to_signed(1, 8),
    to_signed(2, 8),
    to_signed(1, 8),
    to_signed(-1, 8),
    to_signed(-4, 8),
    to_signed(-6, 8),
    to_signed(-7, 8),
    to_signed(-6, 8),
    to_signed(-3, 8),
    to_signed(0, 8),
    to_signed(3, 8),
    to_signed(5, 8),
    to_signed(5, 8),
    to_signed(3, 8),
    to_signed(-1, 8),
    to_signed(-6, 8),
    to_signed(-10, 8),
    to_signed(-12, 8),
    to_signed(-12, 8),
    to_signed(-10, 8),
    to_signed(-6, 8),
    to_signed(-2, 8),
    to_signed(1, 8),
    to_signed(3, 8),
    to_signed(2, 8),
    to_signed(0, 8),
    to_signed(-3, 8),
    to_signed(-5, 8),
    to_signed(-5, 8),
    to_signed(-3, 8),
    to_signed(1, 8),
    to_signed(6, 8),
    to_signed(12, 8),
    to_signed(16, 8),
    to_signed(17, 8),
    to_signed(15, 8),
    to_signed(13, 8),
    to_signed(9, 8),
    to_signed(5, 8),
    to_signed(0, 8),
    to_signed(-2, 8),
    to_signed(-1, 8),
    to_signed(0, 8),
    to_signed(2, 8),
    to_signed(6, 8),
    to_signed(9, 8),
    to_signed(10, 8),
    to_signed(8, 8),
    to_signed(6, 8),
    to_signed(3, 8),
    to_signed(0, 8),
    to_signed(-1, 8),
    to_signed(0, 8),
    to_signed(2, 8),
    to_signed(4, 8),
    to_signed(6, 8),
    to_signed(8, 8),
    to_signed(8, 8),
    to_signed(5, 8),
    to_signed(1, 8),
    to_signed(-1, 8),
    to_signed(-3, 8),
    to_signed(-4, 8),
    to_signed(-4, 8),
    to_signed(-2, 8),
    to_signed(0, 8),
    to_signed(1, 8),
    to_signed(0, 8),
    to_signed(0, 8),
    to_signed(1, 8),
    to_signed(2, 8),
    to_signed(3, 8),
    to_signed(5, 8),
    to_signed(5, 8),
    to_signed(4, 8),
    to_signed(4, 8),
    to_signed(4, 8),
    to_signed(4, 8),
    to_signed(3, 8),
    to_signed(3, 8),
    to_signed(3, 8),
    to_signed(0, 8),
    to_signed(-4, 8),
    to_signed(-7, 8),
    to_signed(-7, 8),
    to_signed(-5, 8),
    to_signed(-4, 8),
    to_signed(-2, 8),
    to_signed(-1, 8),
    to_signed(-2, 8),
    to_signed(-6, 8),
    to_signed(-10, 8),
    to_signed(-12, 8),
    to_signed(-13, 8),
    to_signed(-12, 8),
    to_signed(-10, 8),
    to_signed(-6, 8),
    to_signed(-2, 8),
    to_signed(0, 8),
    to_signed(3, 8),
    to_signed(4, 8),
    to_signed(3, 8),
    to_signed(0, 8),
    to_signed(-4, 8),
    to_signed(-10, 8),
    to_signed(-14, 8),
    to_signed(-13, 8),
    to_signed(-6, 8),
    to_signed(1, 8),
    to_signed(6, 8),
    to_signed(7, 8),
    to_signed(4, 8),
    to_signed(0, 8),
    to_signed(-4, 8),
    to_signed(-8, 8),
    to_signed(-9, 8),
    to_signed(-8, 8),
    to_signed(-6, 8),
    to_signed(-4, 8),
    to_signed(-3, 8),
    to_signed(-3, 8),
    to_signed(-2, 8),
    to_signed(-1, 8),
    to_signed(-1, 8),
    to_signed(-3, 8),
    to_signed(-6, 8),
    to_signed(-9, 8),
    to_signed(-12, 8),
    to_signed(-11, 8),
    to_signed(-7, 8),
    to_signed(-2, 8),
    to_signed(2, 8),
    to_signed(3, 8),
    to_signed(2, 8),
    to_signed(-1, 8),
    to_signed(-5, 8),
    to_signed(-8, 8),
    to_signed(-8, 8),
    to_signed(-7, 8),
    to_signed(-4, 8),
    to_signed(0, 8),
    to_signed(5, 8),
    to_signed(8, 8),
    to_signed(8, 8),
    to_signed(7, 8),
    to_signed(6, 8),
    to_signed(3, 8),
    to_signed(-1, 8),
    to_signed(-4, 8),
    to_signed(-5, 8),
    to_signed(-4, 8),
    to_signed(0, 8),
    to_signed(5, 8),
    to_signed(10, 8),
    to_signed(9, 8),
    to_signed(5, 8),
    to_signed(-1, 8),
    to_signed(-5, 8),
    to_signed(-9, 8),
    to_signed(-12, 8),
    to_signed(-11, 8),
    to_signed(-6, 8),
    to_signed(-2, 8),
    to_signed(1, 8),
    to_signed(3, 8),
    to_signed(2, 8),
    to_signed(-1, 8),
    to_signed(-5, 8),
    to_signed(-7, 8),
    to_signed(-10, 8),
    to_signed(-13, 8),
    to_signed(-14, 8),
    to_signed(-12, 8),
    to_signed(-8, 8),
    to_signed(-5, 8),
    to_signed(-3, 8),
    to_signed(-2, 8),
    to_signed(-3, 8),
    to_signed(-5, 8),
    to_signed(-7, 8),
    to_signed(-9, 8),
    to_signed(-10, 8),
    to_signed(-10, 8),
    to_signed(-7, 8),
    to_signed(-3, 8),
    to_signed(2, 8),
    to_signed(6, 8),
    to_signed(8, 8),
    to_signed(8, 8),
    to_signed(6, 8),
    to_signed(3, 8),
    to_signed(0, 8),
    to_signed(-4, 8),
    to_signed(-6, 8),
    to_signed(-6, 8),
    to_signed(-4, 8),
    to_signed(-2, 8),
    to_signed(1, 8),
    to_signed(2, 8),
    to_signed(3, 8),
    to_signed(2, 8),
    to_signed(0, 8),
    to_signed(-3, 8),
    to_signed(-5, 8),
    to_signed(-6, 8),
    to_signed(-4, 8),
    to_signed(-1, 8),
    to_signed(2, 8),
    to_signed(6, 8),
    to_signed(9, 8),
    to_signed(9, 8),
    to_signed(6, 8),
    to_signed(1, 8),
    to_signed(-4, 8),
    to_signed(-7, 8),
    to_signed(-9, 8),
    to_signed(-8, 8),
    to_signed(-4, 8),
    to_signed(1, 8),
    to_signed(3, 8),
    to_signed(1, 8),
    to_signed(-3, 8),
    to_signed(-8, 8),
    to_signed(-11, 8),
    to_signed(-13, 8),
    to_signed(-14, 8),
    to_signed(-13, 8),
    to_signed(-11, 8),
    to_signed(-9, 8),
    to_signed(-6, 8),
    to_signed(-3, 8),
    to_signed(-2, 8),
    to_signed(-2, 8),
    to_signed(-4, 8),
    to_signed(-8, 8),
    to_signed(-13, 8),
    to_signed(-17, 8),
    to_signed(-18, 8),
    to_signed(-16, 8),
    to_signed(-12, 8),
    to_signed(-7, 8),
    to_signed(-3, 8),
    to_signed(-2, 8),
    to_signed(-4, 8),
    to_signed(-6, 8),
    to_signed(-8, 8),
    to_signed(-11, 8),
    to_signed(-13, 8),
    to_signed(-14, 8),
    to_signed(-12, 8),
    to_signed(-9, 8),
    to_signed(-6, 8),
    to_signed(-1, 8),
    to_signed(3, 8),
    to_signed(5, 8),
    to_signed(4, 8),
    to_signed(1, 8),
    to_signed(-4, 8),
    to_signed(-8, 8),
    to_signed(-10, 8),
    to_signed(-7, 8),
    to_signed(-2, 8),
    to_signed(5, 8),
    to_signed(11, 8),
    to_signed(13, 8),
    to_signed(12, 8),
    to_signed(8, 8),
    to_signed(4, 8),
    to_signed(2, 8),
    to_signed(1, 8),
    to_signed(1, 8),
    to_signed(3, 8),
    to_signed(5, 8),
    to_signed(7, 8),
    to_signed(9, 8),
    to_signed(11, 8),
    to_signed(12, 8),
    to_signed(11, 8),
    to_signed(10, 8),
    to_signed(7, 8),
    to_signed(3, 8),
    to_signed(0, 8),
    to_signed(-1, 8),
    to_signed(0, 8),
    to_signed(2, 8),
    to_signed(4, 8),
    to_signed(6, 8),
    to_signed(6, 8),
    to_signed(4, 8),
    to_signed(1, 8),
    to_signed(-1, 8),
    to_signed(-3, 8),
    to_signed(-4, 8),
    to_signed(-3, 8),
    to_signed(0, 8),
    to_signed(2, 8),
    to_signed(4, 8),
    to_signed(4, 8),
    to_signed(5, 8),
    to_signed(4, 8),
    to_signed(3, 8),
    to_signed(3, 8),
    to_signed(3, 8),
    to_signed(2, 8),
    to_signed(2, 8),
    to_signed(4, 8),
    to_signed(9, 8),
    to_signed(13, 8),
    to_signed(14, 8),
    to_signed(12, 8),
    to_signed(9, 8),
    to_signed(4, 8),
    to_signed(-1, 8),
    to_signed(-4, 8),
    to_signed(-4, 8),
    to_signed(0, 8),
    to_signed(6, 8),
    to_signed(10, 8),
    to_signed(12, 8),
    to_signed(12, 8),
    to_signed(11, 8),
    to_signed(9, 8),
    to_signed(5, 8),
    to_signed(2, 8),
    to_signed(0, 8),
    to_signed(-1, 8),
    to_signed(0, 8),
    to_signed(3, 8),
    to_signed(6, 8),
    to_signed(9, 8),
    to_signed(12, 8),
    to_signed(12, 8),
    to_signed(9, 8),
    to_signed(5, 8),
    to_signed(1, 8),
    to_signed(-1, 8),
    to_signed(-3, 8),
    to_signed(-2, 8),
    to_signed(3, 8),
    to_signed(9, 8),
    to_signed(13, 8),
    to_signed(15, 8),
    to_signed(14, 8),
    to_signed(12, 8),
    to_signed(7, 8),
    to_signed(1, 8),
    to_signed(-2, 8),
    to_signed(-3, 8),
    to_signed(-3, 8),
    to_signed(-4, 8),
    to_signed(-3, 8),
    to_signed(-1, 8),
    to_signed(2, 8),
    to_signed(2, 8),
    to_signed(0, 8),
    to_signed(-3, 8),
    to_signed(-5, 8),
    to_signed(-7, 8),
    to_signed(-9, 8),
    to_signed(-10, 8),
    to_signed(-8, 8),
    to_signed(-5, 8),
    to_signed(-1, 8),
    to_signed(2, 8),
    to_signed(2, 8),
    to_signed(-1, 8),
    to_signed(-5, 8),
    to_signed(-8, 8),
    to_signed(-10, 8),
    to_signed(-9, 8),
    to_signed(-6, 8),
    to_signed(-3, 8),
    to_signed(0, 8),
    to_signed(0, 8),
    to_signed(0, 8),
    to_signed(-1, 8),
    to_signed(-2, 8),
    to_signed(-2, 8),
    to_signed(-2, 8),
    to_signed(0, 8),
    to_signed(2, 8),
    to_signed(3, 8),
    to_signed(5, 8),
    to_signed(8, 8),
    to_signed(11, 8),
    to_signed(13, 8),
    to_signed(13, 8),
    to_signed(11, 8),
    to_signed(7, 8),
    to_signed(2, 8),
    to_signed(-2, 8),
    to_signed(-3, 8),
    to_signed(-1, 8),
    to_signed(3, 8),
    to_signed(7, 8),
    to_signed(10, 8),
    to_signed(10, 8),
    to_signed(8, 8),
    to_signed(3, 8),
    to_signed(-2, 8),
    to_signed(-5, 8),
    to_signed(-7, 8),
    to_signed(-8, 8),
    to_signed(-8, 8),
    to_signed(-6, 8),
    to_signed(-3, 8),
    to_signed(1, 8),
    to_signed(5, 8),
    to_signed(8, 8),
    to_signed(7, 8),
    to_signed(2, 8),
    to_signed(-5, 8),
    to_signed(-12, 8),
    to_signed(-14, 8),
    to_signed(-11, 8),
    to_signed(-5, 8),
    to_signed(1, 8),
    to_signed(4, 8),
    to_signed(5, 8),
    to_signed(3, 8),
    to_signed(0, 8),
    to_signed(-4, 8),
    to_signed(-7, 8),
    to_signed(-8, 8),
    to_signed(-9, 8),
    to_signed(-10, 8),
    to_signed(-10, 8),
    to_signed(-9, 8),
    to_signed(-6, 8),
    to_signed(-3, 8),
    to_signed(0, 8),
    to_signed(1, 8),
    to_signed(1, 8),
    to_signed(-2, 8),
    to_signed(-5, 8),
    to_signed(-6, 8),
    to_signed(-6, 8),
    to_signed(-4, 8),
    to_signed(-2, 8),
    to_signed(0, 8),
    to_signed(3, 8),
    to_signed(4, 8),
    to_signed(2, 8),
    to_signed(-2, 8),
    to_signed(-4, 8),
    to_signed(-4, 8),
    to_signed(-3, 8),
    to_signed(-2, 8),
    to_signed(0, 8),
    to_signed(3, 8),
    to_signed(6, 8),
    to_signed(7, 8),
    to_signed(7, 8),
    to_signed(8, 8),
    to_signed(9, 8),
    to_signed(9, 8),
    to_signed(6, 8),
    to_signed(3, 8),
    to_signed(3, 8),
    to_signed(4, 8),
    to_signed(6, 8),
    to_signed(7, 8),
    to_signed(7, 8),
    to_signed(6, 8),
    to_signed(2, 8),
    to_signed(-2, 8),
    to_signed(-6, 8),
    to_signed(-9, 8),
    to_signed(-9, 8),
    to_signed(-8, 8),
    to_signed(-7, 8),
    to_signed(-5, 8),
    to_signed(-2, 8),
    to_signed(-2, 8),
    to_signed(-3, 8),
    to_signed(-7, 8),
    to_signed(-11, 8),
    to_signed(-13, 8),
    to_signed(-15, 8),
    to_signed(-14, 8),
    to_signed(-13, 8),
    to_signed(-11, 8),
    to_signed(-9, 8),
    to_signed(-7, 8),
    to_signed(-4, 8),
    to_signed(-2, 8),
    to_signed(-3, 8),
    to_signed(-6, 8),
    to_signed(-10, 8),
    to_signed(-11, 8),
    to_signed(-11, 8),
    to_signed(-9, 8),
    to_signed(-4, 8),
    to_signed(1, 8),
    to_signed(5, 8),
    to_signed(7, 8),
    to_signed(7, 8),
    to_signed(6, 8),
    to_signed(3, 8),
    to_signed(1, 8),
    to_signed(-1, 8),
    to_signed(-2, 8),
    to_signed(-4, 8),
    to_signed(-5, 8),
    to_signed(-3, 8),
    to_signed(-1, 8),
    to_signed(1, 8),
    to_signed(2, 8),
    to_signed(2, 8),
    to_signed(1, 8),
    to_signed(-1, 8),
    to_signed(-3, 8),
    to_signed(-6, 8),
    to_signed(-7, 8),
    to_signed(-6, 8),
    to_signed(-3, 8),
    to_signed(0, 8),
    to_signed(1, 8),
    to_signed(0, 8),
    to_signed(-3, 8),
    to_signed(-6, 8),
    to_signed(-7, 8),
    to_signed(-8, 8),
    to_signed(-8, 8),
    to_signed(-7, 8),
    to_signed(-6, 8),
    to_signed(-6, 8),
    to_signed(-7, 8),
    to_signed(-9, 8),
    to_signed(-9, 8),
    to_signed(-10, 8),
    to_signed(-13, 8),
    to_signed(-15, 8),
    to_signed(-15, 8),
    to_signed(-14, 8),
    to_signed(-12, 8),
    to_signed(-10, 8),
    to_signed(-8, 8),
    to_signed(-7, 8),
    to_signed(-7, 8),
    to_signed(-8, 8),
    to_signed(-10, 8),
    to_signed(-13, 8),
    to_signed(-16, 8),
    to_signed(-17, 8),
    to_signed(-17, 8),
    to_signed(-15, 8),
    to_signed(-11, 8),
    to_signed(-6, 8),
    to_signed(-3, 8),
    to_signed(-3, 8),
    to_signed(-6, 8),
    to_signed(-11, 8),
    to_signed(-14, 8),
    to_signed(-16, 8),
    to_signed(-15, 8),
    to_signed(-12, 8),
    to_signed(-8, 8),
    to_signed(-5, 8),
    to_signed(-2, 8),
    to_signed(2, 8),
    to_signed(7, 8),
    to_signed(9, 8),
    to_signed(8, 8),
    to_signed(6, 8),
    to_signed(4, 8),
    to_signed(4, 8),
    to_signed(5, 8),
    to_signed(8, 8),
    to_signed(13, 8),
    to_signed(20, 8),
    to_signed(26, 8),
    to_signed(28, 8),
    to_signed(27, 8),
    to_signed(24, 8),
    to_signed(21, 8),
    to_signed(17, 8),
    to_signed(13, 8),
    to_signed(12, 8),
    to_signed(12, 8),
    to_signed(13, 8),
    to_signed(15, 8),
    to_signed(19, 8),
    to_signed(23, 8),
    to_signed(24, 8),
    to_signed(23, 8),
    to_signed(21, 8),
    to_signed(17, 8),
    to_signed(14, 8),
    to_signed(13, 8),
    to_signed(16, 8),
    to_signed(20, 8),
    to_signed(23, 8),
    to_signed(25, 8),
    to_signed(26, 8),
    to_signed(24, 8),
    to_signed(20, 8),
    to_signed(16, 8),
    to_signed(14, 8),
    to_signed(14, 8),
    to_signed(14, 8),
    to_signed(14, 8),
    to_signed(15, 8),
    to_signed(17, 8),
    to_signed(18, 8),
    to_signed(19, 8),
    to_signed(19, 8),
    to_signed(18, 8),
    to_signed(16, 8),
    to_signed(15, 8),
    to_signed(17, 8),
    to_signed(18, 8),
    to_signed(17, 8),
    to_signed(18, 8),
    to_signed(20, 8),
    to_signed(21, 8),
    to_signed(20, 8),
    to_signed(18, 8),
    to_signed(15, 8),
    to_signed(10, 8),
    to_signed(3, 8),
    to_signed(-3, 8),
    to_signed(-4, 8),
    to_signed(-2, 8),
    to_signed(2, 8),
    to_signed(5, 8),
    to_signed(5, 8),
    to_signed(2, 8),
    to_signed(-3, 8),
    to_signed(-6, 8),
    to_signed(-9, 8),
    to_signed(-13, 8),
    to_signed(-18, 8),
    to_signed(-20, 8),
    to_signed(-19, 8),
    to_signed(-17, 8),
    to_signed(-13, 8),
    to_signed(-9, 8),
    to_signed(-8, 8),
    to_signed(-9, 8),
    to_signed(-13, 8),
    to_signed(-18, 8),
    to_signed(-23, 8),
    to_signed(-25, 8),
    to_signed(-24, 8),
    to_signed(-22, 8),
    to_signed(-18, 8),
    to_signed(-14, 8),
    to_signed(-12, 8),
    to_signed(-10, 8),
    to_signed(-9, 8),
    to_signed(-10, 8),
    to_signed(-13, 8),
    to_signed(-17, 8),
    to_signed(-19, 8),
    to_signed(-19, 8),
    to_signed(-18, 8),
    to_signed(-17, 8),
    to_signed(-15, 8),
    to_signed(-13, 8),
    to_signed(-9, 8),
    to_signed(-7, 8),
    to_signed(-6, 8),
    to_signed(-6, 8),
    to_signed(-7, 8),
    to_signed(-10, 8),
    to_signed(-12, 8),
    to_signed(-12, 8),
    to_signed(-8, 8),
    to_signed(-4, 8),
    to_signed(0, 8),
    to_signed(2, 8),
    to_signed(3, 8),
    to_signed(2, 8),
    to_signed(1, 8),
    to_signed(1, 8),
    to_signed(0, 8),
    to_signed(0, 8),
    to_signed(2, 8),
    to_signed(6, 8),
    to_signed(8, 8),
    to_signed(7, 8),
    to_signed(6, 8),
    to_signed(5, 8),
    to_signed(4, 8),
    to_signed(1, 8),
    to_signed(-1, 8),
    to_signed(0, 8),
    to_signed(3, 8),
    to_signed(5, 8),
    to_signed(7, 8),
    to_signed(9, 8),
    to_signed(10, 8),
    to_signed(8, 8),
    to_signed(5, 8),
    to_signed(1, 8),
    to_signed(-3, 8),
    to_signed(-7, 8),
    to_signed(-8, 8),
    to_signed(-7, 8),
    to_signed(-4, 8),
    to_signed(-2, 8),
    to_signed(-2, 8),
    to_signed(-3, 8),
    to_signed(-5, 8),
    to_signed(-8, 8),
    to_signed(-13, 8),
    to_signed(-17, 8),
    to_signed(-20, 8),
    to_signed(-21, 8),
    to_signed(-21, 8),
    to_signed(-19, 8),
    to_signed(-16, 8),
    to_signed(-11, 8),
    to_signed(-7, 8),
    to_signed(-4, 8),
    to_signed(-3, 8),
    to_signed(-4, 8),
    to_signed(-6, 8),
    to_signed(-10, 8),
    to_signed(-12, 8),
    to_signed(-10, 8),
    to_signed(-5, 8),
    to_signed(1, 8),
    to_signed(6, 8),
    to_signed(10, 8),
    to_signed(10, 8),
    to_signed(7, 8),
    to_signed(4, 8),
    to_signed(1, 8),
    to_signed(0, 8),
    to_signed(0, 8),
    to_signed(1, 8),
    to_signed(2, 8),
    to_signed(2, 8),
    to_signed(3, 8),
    to_signed(5, 8),
    to_signed(8, 8),
    to_signed(10, 8),
    to_signed(11, 8),
    to_signed(10, 8),
    to_signed(7, 8),
    to_signed(4, 8),
    to_signed(2, 8),
    to_signed(3, 8),
    to_signed(6, 8),
    to_signed(8, 8),
    to_signed(9, 8),
    to_signed(9, 8),
    to_signed(8, 8),
    to_signed(3, 8),
    to_signed(-2, 8),
    to_signed(-4, 8),
    to_signed(-4, 8),
    to_signed(-3, 8),
    to_signed(-1, 8),
    to_signed(1, 8),
    to_signed(2, 8),
    to_signed(1, 8),
    to_signed(0, 8),
    to_signed(-1, 8),
    to_signed(-2, 8),
    to_signed(-5, 8),
    to_signed(-7, 8),
    to_signed(-7, 8),
    to_signed(-5, 8),
    to_signed(-2, 8),
    to_signed(1, 8),
    to_signed(4, 8),
    to_signed(5, 8),
    to_signed(2, 8),
    to_signed(-3, 8),
    to_signed(-8, 8),
    to_signed(-13, 8),
    to_signed(-16, 8),
    to_signed(-16, 8),
    to_signed(-13, 8),
    to_signed(-9, 8),
    to_signed(-5, 8),
    to_signed(-2, 8),
    to_signed(0, 8),
    to_signed(0, 8),
    to_signed(-4, 8),
    to_signed(-11, 8),
    to_signed(-17, 8),
    to_signed(-20, 8),
    to_signed(-20, 8),
    to_signed(-18, 8),
    to_signed(-14, 8),
    to_signed(-8, 8),
    to_signed(-1, 8),
    to_signed(4, 8),
    to_signed(6, 8),
    to_signed(5, 8),
    to_signed(2, 8),
    to_signed(-5, 8),
    to_signed(-11, 8),
    to_signed(-14, 8),
    to_signed(-12, 8),
    to_signed(-5, 8),
    to_signed(3, 8),
    to_signed(9, 8),
    to_signed(11, 8),
    to_signed(11, 8),
    to_signed(8, 8),
    to_signed(6, 8),
    to_signed(4, 8),
    to_signed(2, 8),
    to_signed(-2, 8),
    to_signed(-5, 8),
    to_signed(-6, 8),
    to_signed(-4, 8),
    to_signed(-1, 8),
    to_signed(3, 8),
    to_signed(6, 8),
    to_signed(7, 8),
    to_signed(6, 8),
    to_signed(2, 8),
    to_signed(-3, 8),
    to_signed(-7, 8),
    to_signed(-8, 8),
    to_signed(-6, 8),
    to_signed(-3, 8),
    to_signed(0, 8),
    to_signed(2, 8),
    to_signed(3, 8),
    to_signed(2, 8),
    to_signed(-1, 8),
    to_signed(-4, 8),
    to_signed(-5, 8),
    to_signed(-5, 8),
    to_signed(-3, 8),
    to_signed(0, 8),
    to_signed(3, 8),
    to_signed(5, 8),
    to_signed(5, 8),
    to_signed(5, 8),
    to_signed(4, 8),
    to_signed(3, 8),
    to_signed(1, 8),
    to_signed(-2, 8),
    to_signed(-4, 8),
    to_signed(-2, 8),
    to_signed(1, 8),
    to_signed(4, 8),
    to_signed(6, 8),
    to_signed(5, 8),
    to_signed(2, 8),
    to_signed(-1, 8),
    to_signed(-3, 8),
    to_signed(-5, 8),
    to_signed(-6, 8),
    to_signed(-6, 8),
    to_signed(-6, 8),
    to_signed(-4, 8),
    to_signed(-1, 8),
    to_signed(3, 8),
    to_signed(4, 8),
    to_signed(2, 8),
    to_signed(-2, 8),
    to_signed(-6, 8),
    to_signed(-9, 8),
    to_signed(-11, 8),
    to_signed(-11, 8),
    to_signed(-10, 8),
    to_signed(-7, 8),
    to_signed(-3, 8),
    to_signed(3, 8),
    to_signed(9, 8),
    to_signed(12, 8),
    to_signed(11, 8),
    to_signed(6, 8),
    to_signed(-2, 8),
    to_signed(-8, 8),
    to_signed(-9, 8),
    to_signed(-4, 8),
    to_signed(3, 8),
    to_signed(10, 8),
    to_signed(15, 8),
    to_signed(17, 8),
    to_signed(17, 8),
    to_signed(13, 8),
    to_signed(9, 8),
    to_signed(6, 8),
    to_signed(3, 8),
    to_signed(0, 8),
    to_signed(-2, 8),
    to_signed(0, 8),
    to_signed(3, 8),
    to_signed(8, 8),
    to_signed(13, 8),
    to_signed(16, 8),
    to_signed(14, 8),
    to_signed(9, 8),
    to_signed(3, 8),
    to_signed(-2, 8),
    to_signed(-3, 8),
    to_signed(-2, 8),
    to_signed(1, 8),
    to_signed(5, 8),
    to_signed(9, 8),
    to_signed(10, 8),
    to_signed(9, 8),
    to_signed(4, 8),
    to_signed(0, 8),
    to_signed(-3, 8),
    to_signed(-2, 8),
    to_signed(-1, 8),
    to_signed(-1, 8),
    to_signed(0, 8),
    to_signed(3, 8),
    to_signed(6, 8),
    to_signed(7, 8),
    to_signed(6, 8),
    to_signed(4, 8),
    to_signed(2, 8),
    to_signed(1, 8),
    to_signed(1, 8),
    to_signed(3, 8),
    to_signed(4, 8),
    to_signed(7, 8),
    to_signed(9, 8),
    to_signed(9, 8),
    to_signed(7, 8),
    to_signed(5, 8),
    to_signed(3, 8),
    to_signed(0, 8),
    to_signed(-4, 8),
    to_signed(-7, 8),
    to_signed(-7, 8),
    to_signed(-4, 8),
    to_signed(1, 8),
    to_signed(5, 8),
    to_signed(8, 8),
    to_signed(7, 8),
    to_signed(5, 8),
    to_signed(2, 8),
    to_signed(0, 8),
    to_signed(-1, 8),
    to_signed(-3, 8),
    to_signed(-3, 8),
    to_signed(0, 8),
    to_signed(5, 8),
    to_signed(12, 8),
    to_signed(18, 8),
    to_signed(23, 8),
    to_signed(24, 8),
    to_signed(19, 8),
    to_signed(10, 8),
    to_signed(2, 8),
    to_signed(-1, 8),
    to_signed(1, 8),
    to_signed(6, 8),
    to_signed(13, 8),
    to_signed(20, 8),
    to_signed(24, 8),
    to_signed(26, 8),
    to_signed(24, 8),
    to_signed(20, 8),
    to_signed(15, 8),
    to_signed(9, 8),
    to_signed(4, 8),
    to_signed(0, 8),
    to_signed(1, 8),
    to_signed(5, 8),
    to_signed(10, 8),
    to_signed(14, 8),
    to_signed(16, 8),
    to_signed(16, 8),
    to_signed(12, 8),
    to_signed(6, 8),
    to_signed(1, 8),
    to_signed(-3, 8),
    to_signed(-6, 8),
    to_signed(-5, 8),
    to_signed(-3, 8),
    to_signed(0, 8),
    to_signed(2, 8),
    to_signed(2, 8),
    to_signed(0, 8),
    to_signed(-3, 8),
    to_signed(-6, 8),
    to_signed(-8, 8),
    to_signed(-9, 8),
    to_signed(-8, 8),
    to_signed(-6, 8),
    to_signed(-4, 8),
    to_signed(-4, 8),
    to_signed(-6, 8),
    to_signed(-6, 8),
    to_signed(-6, 8),
    to_signed(-5, 8),
    to_signed(-6, 8),
    to_signed(-6, 8),
    to_signed(-5, 8),
    to_signed(-4, 8),
    to_signed(-3, 8),
    to_signed(-1, 8),
    to_signed(2, 8),
    to_signed(4, 8),
    to_signed(3, 8),
    to_signed(-1, 8),
    to_signed(-5, 8),
    to_signed(-9, 8),
    to_signed(-11, 8),
    to_signed(-11, 8),
    to_signed(-8, 8),
    to_signed(-4, 8),
    to_signed(-1, 8),
    to_signed(-1, 8),
    to_signed(-1, 8),
    to_signed(-4, 8),
    to_signed(-7, 8),
    to_signed(-10, 8),
    to_signed(-12, 8),
    to_signed(-14, 8),
    to_signed(-17, 8),
    to_signed(-18, 8),
    to_signed(-15, 8),
    to_signed(-8, 8),
    to_signed(0, 8),
    to_signed(4, 8),
    to_signed(3, 8),
    to_signed(-3, 8),
    to_signed(-10, 8),
    to_signed(-18, 8),
    to_signed(-22, 8),
    to_signed(-22, 8),
    to_signed(-18, 8),
    to_signed(-10, 8),
    to_signed(-3, 8),
    to_signed(3, 8),
    to_signed(4, 8),
    to_signed(1, 8),
    to_signed(-4, 8),
    to_signed(-6, 8),
    to_signed(-8, 8),
    to_signed(-11, 8),
    to_signed(-15, 8),
    to_signed(-17, 8),
    to_signed(-16, 8),
    to_signed(-12, 8),
    to_signed(-5, 8),
    to_signed(0, 8),
    to_signed(2, 8),
    to_signed(1, 8),
    to_signed(-1, 8),
    to_signed(-3, 8),
    to_signed(-7, 8),
    to_signed(-11, 8),
    to_signed(-14, 8),
    to_signed(-13, 8),
    to_signed(-10, 8),
    to_signed(-6, 8),
    to_signed(-5, 8),
    to_signed(-5, 8),
    to_signed(-5, 8),
    to_signed(-5, 8),
    to_signed(-5, 8),
    to_signed(-5, 8),
    to_signed(-5, 8),
    to_signed(-5, 8),
    to_signed(-4, 8),
    to_signed(-4, 8),
    to_signed(-4, 8),
    to_signed(-4, 8),
    to_signed(-3, 8),
    to_signed(0, 8),
    to_signed(3, 8),
    to_signed(4, 8),
    to_signed(3, 8),
    to_signed(1, 8),
    to_signed(2, 8),
    to_signed(6, 8),
    to_signed(9, 8),
    to_signed(11, 8),
    to_signed(8, 8),
    to_signed(3, 8),
    to_signed(-4, 8),
    to_signed(-7, 8),
    to_signed(-6, 8),
    to_signed(-4, 8),
    to_signed(-3, 8),
    to_signed(-2, 8),
    to_signed(-2, 8),
    to_signed(-1, 8),
    to_signed(-1, 8),
    to_signed(-1, 8),
    to_signed(-1, 8),
    to_signed(-1, 8),
    to_signed(-4, 8),
    to_signed(-7, 8),
    to_signed(-9, 8),
    to_signed(-8, 8),
    to_signed(-6, 8),
    to_signed(-2, 8),
    to_signed(2, 8),
    to_signed(6, 8),
    to_signed(7, 8),
    to_signed(6, 8),
    to_signed(4, 8),
    to_signed(-1, 8),
    to_signed(-6, 8),
    to_signed(-9, 8),
    to_signed(-8, 8),
    to_signed(-5, 8),
    to_signed(-1, 8),
    to_signed(3, 8),
    to_signed(6, 8),
    to_signed(8, 8),
    to_signed(8, 8),
    to_signed(7, 8),
    to_signed(5, 8),
    to_signed(2, 8),
    to_signed(-2, 8),
    to_signed(-5, 8),
    to_signed(-4, 8),
    to_signed(-1, 8),
    to_signed(3, 8),
    to_signed(7, 8),
    to_signed(11, 8),
    to_signed(13, 8),
    to_signed(12, 8),
    to_signed(8, 8),
    to_signed(4, 8),
    to_signed(0, 8),
    to_signed(-3, 8),
    to_signed(-6, 8),
    to_signed(-8, 8),
    to_signed(-6, 8),
    to_signed(-3, 8),
    to_signed(0, 8),
    to_signed(2, 8),
    to_signed(3, 8),
    to_signed(3, 8),
    to_signed(3, 8),
    to_signed(3, 8),
    to_signed(5, 8),
    to_signed(5, 8),
    to_signed(3, 8),
    to_signed(1, 8),
    to_signed(1, 8),
    to_signed(4, 8),
    to_signed(8, 8),
    to_signed(11, 8),
    to_signed(12, 8),
    to_signed(10, 8),
    to_signed(8, 8),
    to_signed(6, 8),
    to_signed(7, 8),
    to_signed(9, 8),
    to_signed(13, 8),
    to_signed(17, 8),
    to_signed(19, 8),
    to_signed(15, 8),
    to_signed(6, 8),
    to_signed(-4, 8),
    to_signed(-9, 8),
    to_signed(-8, 8),
    to_signed(-3, 8),
    to_signed(5, 8),
    to_signed(12, 8),
    to_signed(14, 8),
    to_signed(11, 8),
    to_signed(4, 8),
    to_signed(-3, 8),
    to_signed(-10, 8),
    to_signed(-16, 8),
    to_signed(-17, 8),
    to_signed(-14, 8),
    to_signed(-10, 8),
    to_signed(-5, 8),
    to_signed(-1, 8),
    to_signed(4, 8),
    to_signed(8, 8),
    to_signed(8, 8),
    to_signed(5, 8),
    to_signed(0, 8),
    to_signed(-5, 8),
    to_signed(-7, 8),
    to_signed(-5, 8),
    to_signed(0, 8),
    to_signed(5, 8),
    to_signed(9, 8),
    to_signed(10, 8),
    to_signed(8, 8),
    to_signed(7, 8),
    to_signed(8, 8),
    to_signed(8, 8),
    to_signed(6, 8),
    to_signed(3, 8),
    to_signed(0, 8),
    to_signed(-2, 8),
    to_signed(-4, 8),
    to_signed(-5, 8),
    to_signed(-3, 8),
    to_signed(0, 8),
    to_signed(4, 8),
    to_signed(7, 8),
    to_signed(6, 8),
    to_signed(1, 8),
    to_signed(-4, 8),
    to_signed(-5, 8),
    to_signed(-5, 8),
    to_signed(-5, 8),
    to_signed(-5, 8),
    to_signed(-3, 8),
    to_signed(0, 8),
    to_signed(3, 8),
    to_signed(4, 8),
    to_signed(3, 8),
    to_signed(2, 8),
    to_signed(1, 8),
    to_signed(1, 8),
    to_signed(1, 8),
    to_signed(-2, 8),
    to_signed(-6, 8),
    to_signed(-9, 8),
    to_signed(-7, 8),
    to_signed(-2, 8),
    to_signed(1, 8),
    to_signed(4, 8),
    to_signed(6, 8),
    to_signed(7, 8),
    to_signed(8, 8),
    to_signed(9, 8),
    to_signed(9, 8),
    to_signed(7, 8),
    to_signed(5, 8),
    to_signed(2, 8),
    to_signed(-2, 8),
    to_signed(-6, 8),
    to_signed(-9, 8),
    to_signed(-11, 8),
    to_signed(-11, 8),
    to_signed(-10, 8),
    to_signed(-9, 8),
    to_signed(-8, 8),
    to_signed(-6, 8),
    to_signed(-4, 8),
    to_signed(-3, 8),
    to_signed(-5, 8),
    to_signed(-11, 8),
    to_signed(-19, 8),
    to_signed(-26, 8),
    to_signed(-28, 8),
    to_signed(-27, 8),
    to_signed(-21, 8),
    to_signed(-15, 8),
    to_signed(-11, 8),
    to_signed(-6, 8),
    to_signed(-1, 8),
    to_signed(2, 8),
    to_signed(0, 8),
    to_signed(-6, 8),
    to_signed(-13, 8),
    to_signed(-15, 8),
    to_signed(-14, 8),
    to_signed(-10, 8),
    to_signed(-5, 8),
    to_signed(1, 8),
    to_signed(6, 8),
    to_signed(8, 8),
    to_signed(6, 8),
    to_signed(3, 8),
    to_signed(0, 8),
    to_signed(-2, 8),
    to_signed(-3, 8),
    to_signed(-3, 8),
    to_signed(-4, 8),
    to_signed(-6, 8),
    to_signed(-5, 8),
    to_signed(-3, 8),
    to_signed(1, 8),
    to_signed(4, 8),
    to_signed(7, 8),
    to_signed(8, 8),
    to_signed(6, 8),
    to_signed(3, 8),
    to_signed(1, 8),
    to_signed(-2, 8),
    to_signed(-5, 8),
    to_signed(-7, 8),
    to_signed(-5, 8),
    to_signed(-3, 8),
    to_signed(1, 8),
    to_signed(6, 8),
    to_signed(10, 8),
    to_signed(11, 8),
    to_signed(10, 8),
    to_signed(9, 8),
    to_signed(7, 8),
    to_signed(4, 8),
    to_signed(-1, 8),
    to_signed(-5, 8),
    to_signed(-5, 8),
    to_signed(-2, 8),
    to_signed(3, 8),
    to_signed(5, 8),
    to_signed(6, 8),
    to_signed(5, 8),
    to_signed(3, 8),
    to_signed(1, 8),
    to_signed(0, 8),
    to_signed(0, 8),
    to_signed(3, 8),
    to_signed(4, 8),
    to_signed(2, 8),
    to_signed(-2, 8),
    to_signed(-8, 8),
    to_signed(-13, 8),
    to_signed(-15, 8),
    to_signed(-14, 8),
    to_signed(-10, 8),
    to_signed(-6, 8),
    to_signed(-4, 8),
    to_signed(-3, 8),
    to_signed(-4, 8),
    to_signed(-7, 8),
    to_signed(-14, 8),
    to_signed(-21, 8),
    to_signed(-26, 8),
    to_signed(-28, 8),
    to_signed(-27, 8),
    to_signed(-23, 8),
    to_signed(-20, 8),
    to_signed(-16, 8),
    to_signed(-11, 8),
    to_signed(-6, 8),
    to_signed(-2, 8),
    to_signed(-1, 8),
    to_signed(-4, 8),
    to_signed(-7, 8),
    to_signed(-8, 8),
    to_signed(-7, 8),
    to_signed(-3, 8),
    to_signed(1, 8),
    to_signed(4, 8),
    to_signed(6, 8),
    to_signed(9, 8),
    to_signed(12, 8),
    to_signed(13, 8),
    to_signed(12, 8),
    to_signed(10, 8),
    to_signed(7, 8),
    to_signed(5, 8),
    to_signed(2, 8),
    to_signed(1, 8),
    to_signed(2, 8),
    to_signed(7, 8),
    to_signed(12, 8),
    to_signed(17, 8),
    to_signed(18, 8),
    to_signed(15, 8),
    to_signed(10, 8),
    to_signed(6, 8),
    to_signed(1, 8),
    to_signed(-5, 8),
    to_signed(-11, 8),
    to_signed(-12, 8),
    to_signed(-9, 8),
    to_signed(-3, 8),
    to_signed(5, 8),
    to_signed(10, 8),
    to_signed(12, 8),
    to_signed(10, 8),
    to_signed(6, 8),
    to_signed(2, 8),
    to_signed(-5, 8),
    to_signed(-12, 8),
    to_signed(-18, 8),
    to_signed(-18, 8),
    to_signed(-13, 8),
    to_signed(-4, 8),
    to_signed(5, 8),
    to_signed(10, 8),
    to_signed(9, 8),
    to_signed(6, 8),
    to_signed(3, 8),
    to_signed(1, 8),
    to_signed(2, 8),
    to_signed(5, 8),
    to_signed(7, 8),
    to_signed(4, 8),
    to_signed(-3, 8),
    to_signed(-11, 8),
    to_signed(-18, 8),
    to_signed(-23, 8),
    to_signed(-24, 8),
    to_signed(-21, 8),
    to_signed(-13, 8),
    to_signed(-4, 8),
    to_signed(3, 8),
    to_signed(3, 8),
    to_signed(-3, 8),
    to_signed(-14, 8),
    to_signed(-25, 8),
    to_signed(-33, 8),
    to_signed(-36, 8),
    to_signed(-34, 8),
    to_signed(-26, 8),
    to_signed(-16, 8),
    to_signed(-6, 8),
    to_signed(1, 8),
    to_signed(6, 8),
    to_signed(9, 8),
    to_signed(12, 8),
    to_signed(13, 8),
    to_signed(11, 8),
    to_signed(7, 8),
    to_signed(4, 8),
    to_signed(5, 8),
    to_signed(10, 8),
    to_signed(15, 8),
    to_signed(19, 8),
    to_signed(19, 8),
    to_signed(16, 8),
    to_signed(13, 8),
    to_signed(12, 8),
    to_signed(14, 8),
    to_signed(17, 8),
    to_signed(20, 8),
    to_signed(20, 8),
    to_signed(19, 8),
    to_signed(18, 8),
    to_signed(18, 8),
    to_signed(18, 8),
    to_signed(19, 8),
    to_signed(19, 8),
    to_signed(16, 8),
    to_signed(12, 8),
    to_signed(6, 8),
    to_signed(1, 8),
    to_signed(-4, 8),
    to_signed(-7, 8),
    to_signed(-5, 8),
    to_signed(1, 8),
    to_signed(7, 8),
    to_signed(10, 8),
    to_signed(13, 8),
    to_signed(14, 8),
    to_signed(13, 8),
    to_signed(9, 8),
    to_signed(2, 8),
    to_signed(-7, 8),
    to_signed(-12, 8),
    to_signed(-13, 8),
    to_signed(-7, 8),
    to_signed(2, 8),
    to_signed(11, 8),
    to_signed(22, 8),
    to_signed(30, 8),
    to_signed(33, 8),
    to_signed(32, 8),
    to_signed(27, 8),
    to_signed(20, 8),
    to_signed(14, 8),
    to_signed(11, 8),
    to_signed(10, 8),
    to_signed(7, 8),
    to_signed(0, 8),
    to_signed(-9, 8),
    to_signed(-14, 8),
    to_signed(-14, 8),
    to_signed(-9, 8),
    to_signed(1, 8),
    to_signed(10, 8),
    to_signed(16, 8),
    to_signed(15, 8),
    to_signed(6, 8),
    to_signed(-7, 8),
    to_signed(-21, 8),
    to_signed(-30, 8),
    to_signed(-32, 8),
    to_signed(-28, 8),
    to_signed(-21, 8),
    to_signed(-15, 8),
    to_signed(-10, 8),
    to_signed(-4, 8),
    to_signed(3, 8),
    to_signed(10, 8),
    to_signed(12, 8),
    to_signed(10, 8),
    to_signed(6, 8),
    to_signed(3, 8),
    to_signed(3, 8),
    to_signed(3, 8),
    to_signed(3, 8),
    to_signed(4, 8),
    to_signed(8, 8),
    to_signed(11, 8),
    to_signed(11, 8),
    to_signed(11, 8),
    to_signed(11, 8),
    to_signed(14, 8),
    to_signed(18, 8),
    to_signed(19, 8),
    to_signed(15, 8),
    to_signed(9, 8),
    to_signed(5, 8),
    to_signed(6, 8),
    to_signed(9, 8),
    to_signed(11, 8),
    to_signed(10, 8),
    to_signed(8, 8),
    to_signed(5, 8),
    to_signed(-1, 8),
    to_signed(-9, 8),
    to_signed(-17, 8),
    to_signed(-22, 8),
    to_signed(-19, 8),
    to_signed(-11, 8),
    to_signed(1, 8),
    to_signed(11, 8),
    to_signed(17, 8),
    to_signed(20, 8),
    to_signed(19, 8),
    to_signed(14, 8),
    to_signed(3, 8),
    to_signed(-10, 8),
    to_signed(-20, 8),
    to_signed(-24, 8),
    to_signed(-19, 8),
    to_signed(-8, 8),
    to_signed(3, 8),
    to_signed(10, 8),
    to_signed(14, 8),
    to_signed(16, 8),
    to_signed(17, 8),
    to_signed(16, 8),
    to_signed(14, 8),
    to_signed(11, 8),
    to_signed(6, 8),
    to_signed(-2, 8),
    to_signed(-11, 8),
    to_signed(-20, 8),
    to_signed(-27, 8),
    to_signed(-29, 8),
    to_signed(-25, 8),
    to_signed(-16, 8),
    to_signed(-8, 8),
    to_signed(-2, 8),
    to_signed(1, 8),
    to_signed(-1, 8),
    to_signed(-8, 8),
    to_signed(-20, 8),
    to_signed(-32, 8),
    to_signed(-40, 8),
    to_signed(-41, 8),
    to_signed(-35, 8),
    to_signed(-27, 8),
    to_signed(-20, 8),
    to_signed(-12, 8),
    to_signed(-2, 8),
    to_signed(9, 8),
    to_signed(17, 8),
    to_signed(18, 8),
    to_signed(12, 8),
    to_signed(4, 8),
    to_signed(1, 8),
    to_signed(2, 8),
    to_signed(5, 8),
    to_signed(9, 8),
    to_signed(10, 8),
    to_signed(10, 8),
    to_signed(8, 8),
    to_signed(9, 8),
    to_signed(14, 8),
    to_signed(20, 8),
    to_signed(24, 8),
    to_signed(24, 8),
    to_signed(19, 8),
    to_signed(13, 8),
    to_signed(8, 8),
    to_signed(7, 8),
    to_signed(6, 8),
    to_signed(6, 8),
    to_signed(5, 8),
    to_signed(6, 8),
    to_signed(7, 8),
    to_signed(8, 8),
    to_signed(6, 8),
    to_signed(-1, 8),
    to_signed(-12, 8),
    to_signed(-22, 8),
    to_signed(-25, 8),
    to_signed(-18, 8),
    to_signed(-5, 8),
    to_signed(8, 8),
    to_signed(14, 8),
    to_signed(12, 8),
    to_signed(7, 8),
    to_signed(1, 8),
    to_signed(-4, 8),
    to_signed(-12, 8),
    to_signed(-23, 8),
    to_signed(-31, 8),
    to_signed(-30, 8),
    to_signed(-21, 8),
    to_signed(-8, 8),
    to_signed(2, 8),
    to_signed(7, 8),
    to_signed(9, 8),
    to_signed(10, 8),
    to_signed(10, 8),
    to_signed(10, 8),
    to_signed(6, 8),
    to_signed(2, 8),
    to_signed(-4, 8),
    to_signed(-12, 8),
    to_signed(-21, 8),
    to_signed(-30, 8),
    to_signed(-33, 8),
    to_signed(-30, 8),
    to_signed(-23, 8),
    to_signed(-14, 8),
    to_signed(-8, 8),
    to_signed(-4, 8),
    to_signed(-4, 8),
    to_signed(-8, 8),
    to_signed(-18, 8),
    to_signed(-30, 8),
    to_signed(-40, 8),
    to_signed(-42, 8),
    to_signed(-38, 8),
    to_signed(-31, 8),
    to_signed(-24, 8),
    to_signed(-14, 8),
    to_signed(-4, 8),
    to_signed(7, 8),
    to_signed(14, 8),
    to_signed(16, 8),
    to_signed(15, 8),
    to_signed(12, 8),
    to_signed(10, 8),
    to_signed(9, 8),
    to_signed(10, 8),
    to_signed(12, 8),
    to_signed(12, 8),
    to_signed(11, 8),
    to_signed(9, 8),
    to_signed(6, 8),
    to_signed(5, 8),
    to_signed(6, 8),
    to_signed(10, 8),
    to_signed(15, 8),
    to_signed(21, 8),
    to_signed(24, 8),
    to_signed(23, 8),
    to_signed(18, 8),
    to_signed(11, 8),
    to_signed(7, 8),
    to_signed(7, 8),
    to_signed(9, 8),
    to_signed(9, 8),
    to_signed(4, 8),
    to_signed(-7, 8),
    to_signed(-21, 8),
    to_signed(-33, 8),
    to_signed(-38, 8),
    to_signed(-33, 8),
    to_signed(-20, 8),
    to_signed(-5, 8),
    to_signed(5, 8),
    to_signed(10, 8),
    to_signed(13, 8),
    to_signed(14, 8),
    to_signed(9, 8),
    to_signed(-5, 8),
    to_signed(-24, 8),
    to_signed(-40, 8),
    to_signed(-45, 8),
    to_signed(-38, 8),
    to_signed(-24, 8),
    to_signed(-11, 8),
    to_signed(0, 8),
    to_signed(8, 8),
    to_signed(16, 8),
    to_signed(19, 8),
    to_signed(16, 8),
    to_signed(10, 8),
    to_signed(5, 8),
    to_signed(0, 8),
    to_signed(-7, 8),
    to_signed(-19, 8),
    to_signed(-33, 8),
    to_signed(-43, 8),
    to_signed(-45, 8),
    to_signed(-41, 8),
    to_signed(-33, 8),
    to_signed(-23, 8),
    to_signed(-12, 8),
    to_signed(-4, 8),
    to_signed(-2, 8),
    to_signed(-10, 8),
    to_signed(-22, 8),
    to_signed(-33, 8),
    to_signed(-39, 8),
    to_signed(-40, 8),
    to_signed(-40, 8),
    to_signed(-37, 8),
    to_signed(-29, 8),
    to_signed(-15, 8),
    to_signed(0, 8),
    to_signed(13, 8),
    to_signed(20, 8),
    to_signed(21, 8),
    to_signed(21, 8),
    to_signed(22, 8),
    to_signed(22, 8),
    to_signed(20, 8),
    to_signed(17, 8),
    to_signed(14, 8),
    to_signed(14, 8),
    to_signed(15, 8),
    to_signed(17, 8),
    to_signed(19, 8),
    to_signed(20, 8),
    to_signed(23, 8),
    to_signed(28, 8),
    to_signed(33, 8),
    to_signed(36, 8),
    to_signed(35, 8),
    to_signed(31, 8),
    to_signed(27, 8),
    to_signed(24, 8),
    to_signed(23, 8),
    to_signed(22, 8),
    to_signed(19, 8),
    to_signed(15, 8),
    to_signed(7, 8),
    to_signed(-5, 8),
    to_signed(-19, 8),
    to_signed(-29, 8),
    to_signed(-29, 8),
    to_signed(-17, 8),
    to_signed(0, 8),
    to_signed(15, 8),
    to_signed(26, 8),
    to_signed(34, 8),
    to_signed(39, 8),
    to_signed(38, 8),
    to_signed(27, 8),
    to_signed(7, 8),
    to_signed(-15, 8),
    to_signed(-30, 8),
    to_signed(-33, 8),
    to_signed(-28, 8),
    to_signed(-18, 8),
    to_signed(-6, 8),
    to_signed(9, 8),
    to_signed(22, 8),
    to_signed(31, 8),
    to_signed(32, 8),
    to_signed(28, 8),
    to_signed(22, 8),
    to_signed(15, 8),
    to_signed(5, 8),
    to_signed(-9, 8),
    to_signed(-25, 8),
    to_signed(-37, 8),
    to_signed(-40, 8),
    to_signed(-38, 8),
    to_signed(-34, 8),
    to_signed(-28, 8),
    to_signed(-20, 8),
    to_signed(-12, 8),
    to_signed(-4, 8),
    to_signed(-2, 8),
    to_signed(-7, 8),
    to_signed(-16, 8),
    to_signed(-27, 8),
    to_signed(-33, 8),
    to_signed(-36, 8),
    to_signed(-34, 8),
    to_signed(-27, 8),
    to_signed(-14, 8),
    to_signed(2, 8),
    to_signed(19, 8),
    to_signed(33, 8),
    to_signed(40, 8),
    to_signed(41, 8),
    to_signed(35, 8),
    to_signed(27, 8),
    to_signed(20, 8),
    to_signed(17, 8),
    to_signed(18, 8),
    to_signed(21, 8),
    to_signed(24, 8),
    to_signed(26, 8),
    to_signed(27, 8),
    to_signed(27, 8),
    to_signed(28, 8),
    to_signed(31, 8),
    to_signed(34, 8),
    to_signed(36, 8),
    to_signed(33, 8),
    to_signed(27, 8),
    to_signed(20, 8),
    to_signed(18, 8),
    to_signed(19, 8),
    to_signed(22, 8),
    to_signed(24, 8),
    to_signed(24, 8),
    to_signed(21, 8),
    to_signed(14, 8),
    to_signed(0, 8),
    to_signed(-18, 8),
    to_signed(-34, 8),
    to_signed(-43, 8),
    to_signed(-39, 8),
    to_signed(-24, 8),
    to_signed(-4, 8),
    to_signed(16, 8),
    to_signed(32, 8),
    to_signed(42, 8),
    to_signed(41, 8),
    to_signed(29, 8),
    to_signed(9, 8),
    to_signed(-13, 8),
    to_signed(-31, 8),
    to_signed(-42, 8),
    to_signed(-43, 8),
    to_signed(-36, 8),
    to_signed(-22, 8),
    to_signed(-6, 8),
    to_signed(8, 8),
    to_signed(19, 8),
    to_signed(24, 8),
    to_signed(26, 8),
    to_signed(24, 8),
    to_signed(18, 8),
    to_signed(8, 8),
    to_signed(-6, 8),
    to_signed(-20, 8),
    to_signed(-34, 8),
    to_signed(-43, 8),
    to_signed(-48, 8),
    to_signed(-47, 8),
    to_signed(-42, 8),
    to_signed(-33, 8),
    to_signed(-22, 8),
    to_signed(-12, 8),
    to_signed(-6, 8),
    to_signed(-5, 8),
    to_signed(-9, 8),
    to_signed(-14, 8),
    to_signed(-21, 8),
    to_signed(-26, 8),
    to_signed(-28, 8),
    to_signed(-25, 8),
    to_signed(-18, 8),
    to_signed(-7, 8),
    to_signed(6, 8),
    to_signed(17, 8),
    to_signed(24, 8),
    to_signed(28, 8),
    to_signed(30, 8),
    to_signed(33, 8),
    to_signed(36, 8),
    to_signed(36, 8),
    to_signed(31, 8),
    to_signed(24, 8),
    to_signed(17, 8),
    to_signed(13, 8),
    to_signed(13, 8),
    to_signed(19, 8),
    to_signed(27, 8),
    to_signed(35, 8),
    to_signed(39, 8),
    to_signed(37, 8),
    to_signed(31, 8),
    to_signed(25, 8),
    to_signed(23, 8),
    to_signed(25, 8),
    to_signed(27, 8),
    to_signed(27, 8),
    to_signed(26, 8),
    to_signed(21, 8),
    to_signed(10, 8),
    to_signed(-7, 8),
    to_signed(-30, 8),
    to_signed(-53, 8),
    to_signed(-65, 8),
    to_signed(-62, 8),
    to_signed(-45, 8),
    to_signed(-19, 8),
    to_signed(8, 8),
    to_signed(32, 8),
    to_signed(46, 8),
    to_signed(47, 8),
    to_signed(34, 8),
    to_signed(9, 8),
    to_signed(-20, 8),
    to_signed(-45, 8),
    to_signed(-60, 8),
    to_signed(-63, 8),
    to_signed(-56, 8),
    to_signed(-41, 8),
    to_signed(-22, 8),
    to_signed(-2, 8),
    to_signed(14, 8),
    to_signed(26, 8),
    to_signed(33, 8),
    to_signed(36, 8),
    to_signed(32, 8),
    to_signed(21, 8),
    to_signed(5, 8),
    to_signed(-13, 8),
    to_signed(-29, 8),
    to_signed(-40, 8),
    to_signed(-47, 8),
    to_signed(-50, 8),
    to_signed(-48, 8),
    to_signed(-39, 8),
    to_signed(-23, 8),
    to_signed(-7, 8),
    to_signed(2, 8),
    to_signed(2, 8),
    to_signed(-5, 8),
    to_signed(-16, 8),
    to_signed(-25, 8),
    to_signed(-34, 8),
    to_signed(-40, 8),
    to_signed(-41, 8),
    to_signed(-33, 8),
    to_signed(-17, 8),
    to_signed(3, 8),
    to_signed(22, 8),
    to_signed(34, 8),
    to_signed(40, 8),
    to_signed(39, 8),
    to_signed(36, 8),
    to_signed(31, 8),
    to_signed(27, 8),
    to_signed(22, 8),
    to_signed(18, 8),
    to_signed(15, 8),
    to_signed(13, 8),
    to_signed(13, 8),
    to_signed(17, 8),
    to_signed(25, 8),
    to_signed(32, 8),
    to_signed(37, 8),
    to_signed(37, 8),
    to_signed(36, 8),
    to_signed(35, 8),
    to_signed(36, 8),
    to_signed(38, 8),
    to_signed(37, 8),
    to_signed(30, 8),
    to_signed(20, 8),
    to_signed(8, 8),
    to_signed(-6, 8),
    to_signed(-25, 8),
    to_signed(-48, 8),
    to_signed(-69, 8),
    to_signed(-80, 8),
    to_signed(-73, 8),
    to_signed(-50, 8),
    to_signed(-21, 8),
    to_signed(7, 8),
    to_signed(30, 8),
    to_signed(44, 8),
    to_signed(47, 8),
    to_signed(36, 8),
    to_signed(11, 8),
    to_signed(-21, 8),
    to_signed(-50, 8),
    to_signed(-66, 8),
    to_signed(-69, 8),
    to_signed(-59, 8),
    to_signed(-41, 8),
    to_signed(-17, 8),
    to_signed(8, 8),
    to_signed(28, 8),
    to_signed(41, 8),
    to_signed(46, 8),
    to_signed(47, 8),
    to_signed(43, 8),
    to_signed(32, 8),
    to_signed(14, 8),
    to_signed(-7, 8),
    to_signed(-25, 8),
    to_signed(-39, 8),
    to_signed(-46, 8),
    to_signed(-48, 8),
    to_signed(-44, 8),
    to_signed(-33, 8),
    to_signed(-19, 8),
    to_signed(-5, 8),
    to_signed(1, 8),
    to_signed(-1, 8),
    to_signed(-11, 8),
    to_signed(-24, 8),
    to_signed(-38, 8),
    to_signed(-49, 8),
    to_signed(-54, 8),
    to_signed(-49, 8),
    to_signed(-35, 8),
    to_signed(-14, 8),
    to_signed(8, 8),
    to_signed(27, 8),
    to_signed(40, 8),
    to_signed(45, 8),
    to_signed(45, 8),
    to_signed(40, 8),
    to_signed(34, 8),
    to_signed(27, 8),
    to_signed(19, 8),
    to_signed(11, 8),
    to_signed(5, 8),
    to_signed(3, 8),
    to_signed(4, 8),
    to_signed(8, 8),
    to_signed(15, 8),
    to_signed(24, 8),
    to_signed(36, 8),
    to_signed(46, 8),
    to_signed(52, 8),
    to_signed(51, 8),
    to_signed(45, 8),
    to_signed(37, 8),
    to_signed(28, 8),
    to_signed(18, 8),
    to_signed(8, 8),
    to_signed(-3, 8),
    to_signed(-16, 8),
    to_signed(-34, 8),
    to_signed(-55, 8),
    to_signed(-72, 8),
    to_signed(-75, 8),
    to_signed(-59, 8),
    to_signed(-28, 8),
    to_signed(5, 8),
    to_signed(30, 8),
    to_signed(43, 8),
    to_signed(47, 8),
    to_signed(41, 8),
    to_signed(23, 8),
    to_signed(-6, 8),
    to_signed(-39, 8),
    to_signed(-63, 8),
    to_signed(-71, 8),
    to_signed(-63, 8),
    to_signed(-45, 8),
    to_signed(-22, 8),
    to_signed(0, 8),
    to_signed(18, 8),
    to_signed(32, 8),
    to_signed(38, 8),
    to_signed(39, 8),
    to_signed(35, 8),
    to_signed(27, 8),
    to_signed(14, 8),
    to_signed(-3, 8),
    to_signed(-20, 8),
    to_signed(-35, 8),
    to_signed(-45, 8),
    to_signed(-49, 8),
    to_signed(-48, 8),
    to_signed(-43, 8),
    to_signed(-33, 8),
    to_signed(-19, 8),
    to_signed(-6, 8),
    to_signed(0, 8),
    to_signed(-3, 8),
    to_signed(-16, 8),
    to_signed(-33, 8),
    to_signed(-49, 8),
    to_signed(-55, 8),
    to_signed(-52, 8),
    to_signed(-41, 8),
    to_signed(-24, 8),
    to_signed(-4, 8),
    to_signed(17, 8),
    to_signed(35, 8),
    to_signed(45, 8),
    to_signed(47, 8),
    to_signed(43, 8),
    to_signed(36, 8),
    to_signed(31, 8),
    to_signed(26, 8),
    to_signed(20, 8),
    to_signed(12, 8),
    to_signed(7, 8),
    to_signed(7, 8),
    to_signed(11, 8),
    to_signed(16, 8),
    to_signed(22, 8),
    to_signed(30, 8),
    to_signed(40, 8),
    to_signed(50, 8),
    to_signed(55, 8),
    to_signed(54, 8),
    to_signed(48, 8),
    to_signed(41, 8),
    to_signed(33, 8),
    to_signed(23, 8),
    to_signed(12, 8),
    to_signed(2, 8),
    to_signed(-9, 8),
    to_signed(-24, 8),
    to_signed(-44, 8),
    to_signed(-64, 8),
    to_signed(-72, 8),
    to_signed(-59, 8),
    to_signed(-28, 8),
    to_signed(9, 8),
    to_signed(37, 8),
    to_signed(53, 8),
    to_signed(57, 8),
    to_signed(50, 8),
    to_signed(33, 8),
    to_signed(7, 8),
    to_signed(-23, 8),
    to_signed(-47, 8),
    to_signed(-60, 8),
    to_signed(-60, 8),
    to_signed(-49, 8),
    to_signed(-33, 8),
    to_signed(-15, 8),
    to_signed(5, 8),
    to_signed(22, 8),
    to_signed(34, 8),
    to_signed(40, 8),
    to_signed(40, 8),
    to_signed(35, 8),
    to_signed(23, 8),
    to_signed(8, 8),
    to_signed(-10, 8),
    to_signed(-27, 8),
    to_signed(-40, 8),
    to_signed(-45, 8),
    to_signed(-42, 8),
    to_signed(-34, 8),
    to_signed(-23, 8),
    to_signed(-13, 8),
    to_signed(-4, 8),
    to_signed(1, 8),
    to_signed(0, 8),
    to_signed(-9, 8),
    to_signed(-25, 8),
    to_signed(-42, 8),
    to_signed(-53, 8),
    to_signed(-55, 8),
    to_signed(-46, 8),
    to_signed(-31, 8),
    to_signed(-11, 8),
    to_signed(10, 8),
    to_signed(29, 8),
    to_signed(41, 8),
    to_signed(45, 8),
    to_signed(43, 8),
    to_signed(39, 8),
    to_signed(34, 8),
    to_signed(28, 8),
    to_signed(21, 8),
    to_signed(14, 8),
    to_signed(11, 8),
    to_signed(14, 8),
    to_signed(19, 8),
    to_signed(24, 8),
    to_signed(30, 8),
    to_signed(36, 8),
    to_signed(46, 8),
    to_signed(55, 8),
    to_signed(61, 8),
    to_signed(63, 8),
    to_signed(61, 8),
    to_signed(56, 8),
    to_signed(48, 8),
    to_signed(36, 8),
    to_signed(21, 8),
    to_signed(2, 8),
    to_signed(-21, 8),
    to_signed(-47, 8),
    to_signed(-71, 8),
    to_signed(-84, 8),
    to_signed(-77, 8),
    to_signed(-52, 8),
    to_signed(-19, 8),
    to_signed(12, 8),
    to_signed(33, 8),
    to_signed(44, 8),
    to_signed(44, 8),
    to_signed(33, 8),
    to_signed(9, 8),
    to_signed(-22, 8),
    to_signed(-50, 8),
    to_signed(-66, 8),
    to_signed(-67, 8),
    to_signed(-55, 8),
    to_signed(-36, 8),
    to_signed(-14, 8),
    to_signed(9, 8),
    to_signed(28, 8),
    to_signed(41, 8),
    to_signed(46, 8),
    to_signed(46, 8),
    to_signed(39, 8),
    to_signed(27, 8),
    to_signed(10, 8),
    to_signed(-10, 8),
    to_signed(-28, 8),
    to_signed(-40, 8),
    to_signed(-44, 8),
    to_signed(-44, 8),
    to_signed(-38, 8),
    to_signed(-29, 8),
    to_signed(-16, 8),
    to_signed(-6, 8),
    to_signed(-3, 8),
    to_signed(-10, 8),
    to_signed(-25, 8),
    to_signed(-43, 8),
    to_signed(-58, 8),
    to_signed(-68, 8),
    to_signed(-69, 8),
    to_signed(-62, 8),
    to_signed(-46, 8),
    to_signed(-23, 8),
    to_signed(2, 8),
    to_signed(27, 8),
    to_signed(44, 8),
    to_signed(53, 8),
    to_signed(54, 8),
    to_signed(49, 8),
    to_signed(43, 8),
    to_signed(37, 8),
    to_signed(30, 8),
    to_signed(24, 8),
    to_signed(19, 8),
    to_signed(16, 8),
    to_signed(17, 8),
    to_signed(20, 8),
    to_signed(24, 8),
    to_signed(31, 8),
    to_signed(40, 8),
    to_signed(49, 8),
    to_signed(56, 8),
    to_signed(57, 8),
    to_signed(54, 8),
    to_signed(50, 8),
    to_signed(45, 8),
    to_signed(38, 8),
    to_signed(28, 8),
    to_signed(14, 8),
    to_signed(-2, 8),
    to_signed(-24, 8),
    to_signed(-50, 8),
    to_signed(-77, 8),
    to_signed(-93, 8),
    to_signed(-88, 8),
    to_signed(-63, 8),
    to_signed(-29, 8),
    to_signed(2, 8),
    to_signed(26, 8),
    to_signed(42, 8),
    to_signed(48, 8),
    to_signed(40, 8),
    to_signed(16, 8),
    to_signed(-18, 8),
    to_signed(-51, 8),
    to_signed(-71, 8),
    to_signed(-75, 8),
    to_signed(-67, 8),
    to_signed(-51, 8),
    to_signed(-30, 8),
    to_signed(-5, 8),
    to_signed(16, 8),
    to_signed(29, 8),
    to_signed(32, 8),
    to_signed(29, 8),
    to_signed(24, 8),
    to_signed(15, 8),
    to_signed(0, 8),
    to_signed(-20, 8),
    to_signed(-41, 8),
    to_signed(-55, 8),
    to_signed(-61, 8),
    to_signed(-60, 8),
    to_signed(-53, 8),
    to_signed(-43, 8),
    to_signed(-29, 8),
    to_signed(-16, 8),
    to_signed(-9, 8),
    to_signed(-9, 8),
    to_signed(-18, 8),
    to_signed(-31, 8),
    to_signed(-44, 8),
    to_signed(-55, 8),
    to_signed(-60, 8),
    to_signed(-58, 8),
    to_signed(-48, 8),
    to_signed(-31, 8),
    to_signed(-8, 8),
    to_signed(16, 8),
    to_signed(38, 8),
    to_signed(54, 8),
    to_signed(61, 8),
    to_signed(61, 8),
    to_signed(56, 8),
    to_signed(49, 8),
    to_signed(39, 8),
    to_signed(28, 8),
    to_signed(18, 8),
    to_signed(12, 8),
    to_signed(11, 8),
    to_signed(13, 8),
    to_signed(18, 8),
    to_signed(24, 8),
    to_signed(33, 8),
    to_signed(44, 8),
    to_signed(52, 8),
    to_signed(54, 8),
    to_signed(53, 8),
    to_signed(50, 8),
    to_signed(49, 8),
    to_signed(45, 8),
    to_signed(38, 8),
    to_signed(26, 8),
    to_signed(9, 8),
    to_signed(-12, 8),
    to_signed(-38, 8),
    to_signed(-66, 8),
    to_signed(-87, 8),
    to_signed(-90, 8),
    to_signed(-73, 8),
    to_signed(-43, 8),
    to_signed(-12, 8),
    to_signed(14, 8),
    to_signed(34, 8),
    to_signed(47, 8),
    to_signed(48, 8),
    to_signed(33, 8),
    to_signed(3, 8),
    to_signed(-32, 8),
    to_signed(-60, 8),
    to_signed(-73, 8),
    to_signed(-74, 8),
    to_signed(-65, 8),
    to_signed(-48, 8),
    to_signed(-26, 8),
    to_signed(-1, 8),
    to_signed(20, 8),
    to_signed(34, 8),
    to_signed(41, 8),
    to_signed(42, 8),
    to_signed(37, 8),
    to_signed(24, 8),
    to_signed(5, 8),
    to_signed(-19, 8),
    to_signed(-41, 8),
    to_signed(-54, 8),
    to_signed(-57, 8),
    to_signed(-50, 8),
    to_signed(-37, 8),
    to_signed(-20, 8),
    to_signed(-3, 8),
    to_signed(9, 8),
    to_signed(13, 8),
    to_signed(8, 8),
    to_signed(-5, 8),
    to_signed(-22, 8),
    to_signed(-39, 8),
    to_signed(-52, 8),
    to_signed(-60, 8),
    to_signed(-61, 8),
    to_signed(-52, 8),
    to_signed(-34, 8),
    to_signed(-6, 8),
    to_signed(23, 8),
    to_signed(46, 8),
    to_signed(58, 8),
    to_signed(59, 8),
    to_signed(56, 8),
    to_signed(53, 8),
    to_signed(46, 8),
    to_signed(34, 8),
    to_signed(19, 8),
    to_signed(7, 8),
    to_signed(1, 8),
    to_signed(3, 8),
    to_signed(10, 8),
    to_signed(18, 8),
    to_signed(29, 8),
    to_signed(42, 8),
    to_signed(53, 8),
    to_signed(58, 8),
    to_signed(57, 8),
    to_signed(53, 8),
    to_signed(50, 8),
    to_signed(48, 8),
    to_signed(42, 8),
    to_signed(29, 8),
    to_signed(11, 8),
    to_signed(-8, 8),
    to_signed(-30, 8),
    to_signed(-54, 8),
    to_signed(-76, 8),
    to_signed(-87, 8),
    to_signed(-80, 8),
    to_signed(-57, 8),
    to_signed(-26, 8),
    to_signed(1, 8),
    to_signed(22, 8),
    to_signed(35, 8),
    to_signed(39, 8),
    to_signed(30, 8),
    to_signed(7, 8),
    to_signed(-23, 8),
    to_signed(-50, 8),
    to_signed(-63, 8),
    to_signed(-62, 8),
    to_signed(-54, 8),
    to_signed(-42, 8),
    to_signed(-26, 8),
    to_signed(-6, 8),
    to_signed(17, 8),
    to_signed(36, 8),
    to_signed(47, 8),
    to_signed(50, 8),
    to_signed(47, 8),
    to_signed(38, 8),
    to_signed(24, 8),
    to_signed(4, 8),
    to_signed(-18, 8),
    to_signed(-36, 8),
    to_signed(-45, 8),
    to_signed(-44, 8),
    to_signed(-35, 8),
    to_signed(-22, 8),
    to_signed(-9, 8),
    to_signed(3, 8),
    to_signed(11, 8),
    to_signed(10, 8),
    to_signed(1, 8),
    to_signed(-16, 8),
    to_signed(-32, 8),
    to_signed(-44, 8),
    to_signed(-50, 8),
    to_signed(-51, 8),
    to_signed(-44, 8),
    to_signed(-29, 8),
    to_signed(-5, 8),
    to_signed(25, 8),
    to_signed(50, 8),
    to_signed(63, 8),
    to_signed(65, 8),
    to_signed(61, 8),
    to_signed(56, 8),
    to_signed(49, 8),
    to_signed(37, 8),
    to_signed(22, 8),
    to_signed(8, 8),
    to_signed(-1, 8),
    to_signed(-3, 8),
    to_signed(0, 8),
    to_signed(6, 8),
    to_signed(16, 8),
    to_signed(30, 8),
    to_signed(45, 8),
    to_signed(55, 8),
    to_signed(58, 8),
    to_signed(57, 8),
    to_signed(55, 8),
    to_signed(51, 8),
    to_signed(40, 8),
    to_signed(22, 8),
    to_signed(1, 8),
    to_signed(-18, 8),
    to_signed(-37, 8),
    to_signed(-56, 8),
    to_signed(-76, 8),
    to_signed(-89, 8),
    to_signed(-85, 8),
    to_signed(-64, 8),
    to_signed(-33, 8),
    to_signed(-4, 8),
    to_signed(17, 8),
    to_signed(30, 8),
    to_signed(34, 8),
    to_signed(27, 8),
    to_signed(9, 8),
    to_signed(-17, 8),
    to_signed(-40, 8),
    to_signed(-54, 8),
    to_signed(-56, 8),
    to_signed(-50, 8),
    to_signed(-39, 8),
    to_signed(-24, 8),
    to_signed(-7, 8),
    to_signed(12, 8),
    to_signed(27, 8),
    to_signed(34, 8),
    to_signed(34, 8),
    to_signed(29, 8),
    to_signed(21, 8),
    to_signed(9, 8),
    to_signed(-7, 8),
    to_signed(-24, 8),
    to_signed(-37, 8),
    to_signed(-43, 8),
    to_signed(-40, 8),
    to_signed(-33, 8),
    to_signed(-22, 8),
    to_signed(-11, 8),
    to_signed(0, 8),
    to_signed(8, 8),
    to_signed(9, 8),
    to_signed(1, 8),
    to_signed(-14, 8),
    to_signed(-31, 8),
    to_signed(-43, 8),
    to_signed(-48, 8),
    to_signed(-48, 8),
    to_signed(-41, 8),
    to_signed(-25, 8),
    to_signed(-1, 8),
    to_signed(27, 8),
    to_signed(50, 8),
    to_signed(61, 8),
    to_signed(61, 8),
    to_signed(55, 8),
    to_signed(48, 8),
    to_signed(40, 8),
    to_signed(30, 8),
    to_signed(18, 8),
    to_signed(7, 8),
    to_signed(2, 8),
    to_signed(1, 8),
    to_signed(4, 8),
    to_signed(9, 8),
    to_signed(17, 8),
    to_signed(28, 8),
    to_signed(37, 8),
    to_signed(41, 8),
    to_signed(42, 8),
    to_signed(41, 8),
    to_signed(41, 8),
    to_signed(37, 8),
    to_signed(26, 8),
    to_signed(10, 8),
    to_signed(-7, 8),
    to_signed(-24, 8),
    to_signed(-40, 8),
    to_signed(-59, 8),
    to_signed(-77, 8),
    to_signed(-86, 8),
    to_signed(-77, 8),
    to_signed(-53, 8),
    to_signed(-23, 8),
    to_signed(2, 8),
    to_signed(19, 8),
    to_signed(27, 8),
    to_signed(28, 8),
    to_signed(20, 8),
    to_signed(3, 8),
    to_signed(-19, 8),
    to_signed(-38, 8),
    to_signed(-47, 8),
    to_signed(-46, 8),
    to_signed(-37, 8),
    to_signed(-26, 8),
    to_signed(-13, 8),
    to_signed(2, 8),
    to_signed(16, 8),
    to_signed(26, 8),
    to_signed(32, 8),
    to_signed(34, 8),
    to_signed(31, 8),
    to_signed(23, 8),
    to_signed(11, 8),
    to_signed(-6, 8),
    to_signed(-22, 8),
    to_signed(-34, 8),
    to_signed(-38, 8),
    to_signed(-34, 8),
    to_signed(-24, 8),
    to_signed(-12, 8),
    to_signed(-1, 8),
    to_signed(8, 8),
    to_signed(12, 8),
    to_signed(8, 8),
    to_signed(-2, 8),
    to_signed(-17, 8),
    to_signed(-32, 8),
    to_signed(-42, 8),
    to_signed(-46, 8),
    to_signed(-43, 8),
    to_signed(-33, 8),
    to_signed(-15, 8),
    to_signed(8, 8),
    to_signed(33, 8),
    to_signed(52, 8),
    to_signed(61, 8),
    to_signed(63, 8),
    to_signed(60, 8),
    to_signed(55, 8),
    to_signed(45, 8),
    to_signed(31, 8),
    to_signed(14, 8),
    to_signed(0, 8),
    to_signed(-7, 8),
    to_signed(-8, 8),
    to_signed(-4, 8),
    to_signed(3, 8),
    to_signed(14, 8),
    to_signed(27, 8),
    to_signed(39, 8),
    to_signed(46, 8),
    to_signed(48, 8),
    to_signed(47, 8),
    to_signed(43, 8),
    to_signed(35, 8),
    to_signed(22, 8),
    to_signed(5, 8),
    to_signed(-11, 8),
    to_signed(-25, 8),
    to_signed(-41, 8),
    to_signed(-58, 8),
    to_signed(-71, 8),
    to_signed(-71, 8),
    to_signed(-54, 8),
    to_signed(-27, 8),
    to_signed(1, 8),
    to_signed(21, 8),
    to_signed(32, 8),
    to_signed(35, 8),
    to_signed(31, 8),
    to_signed(18, 8),
    to_signed(-4, 8),
    to_signed(-29, 8),
    to_signed(-47, 8),
    to_signed(-54, 8),
    to_signed(-48, 8),
    to_signed(-33, 8),
    to_signed(-15, 8),
    to_signed(5, 8),
    to_signed(22, 8),
    to_signed(34, 8),
    to_signed(41, 8),
    to_signed(41, 8),
    to_signed(37, 8),
    to_signed(28, 8),
    to_signed(17, 8),
    to_signed(3, 8),
    to_signed(-10, 8),
    to_signed(-22, 8),
    to_signed(-28, 8),
    to_signed(-28, 8),
    to_signed(-21, 8),
    to_signed(-10, 8),
    to_signed(3, 8),
    to_signed(15, 8),
    to_signed(20, 8),
    to_signed(18, 8),
    to_signed(7, 8),
    to_signed(-8, 8),
    to_signed(-26, 8),
    to_signed(-41, 8),
    to_signed(-50, 8),
    to_signed(-51, 8),
    to_signed(-45, 8),
    to_signed(-31, 8),
    to_signed(-10, 8),
    to_signed(13, 8),
    to_signed(33, 8),
    to_signed(47, 8),
    to_signed(54, 8),
    to_signed(55, 8),
    to_signed(51, 8),
    to_signed(45, 8),
    to_signed(36, 8),
    to_signed(22, 8),
    to_signed(8, 8),
    to_signed(-2, 8),
    to_signed(-6, 8),
    to_signed(-3, 8),
    to_signed(3, 8),
    to_signed(12, 8),
    to_signed(24, 8),
    to_signed(38, 8),
    to_signed(49, 8),
    to_signed(56, 8),
    to_signed(58, 8),
    to_signed(54, 8),
    to_signed(47, 8),
    to_signed(36, 8),
    to_signed(21, 8),
    to_signed(1, 8),
    to_signed(-20, 8),
    to_signed(-42, 8),
    to_signed(-64, 8),
    to_signed(-81, 8),
    to_signed(-87, 8),
    to_signed(-76, 8),
    to_signed(-51, 8),
    to_signed(-21, 8),
    to_signed(5, 8),
    to_signed(22, 8),
    to_signed(28, 8),
    to_signed(26, 8),
    to_signed(16, 8),
    to_signed(-1, 8),
    to_signed(-23, 8),
    to_signed(-43, 8),
    to_signed(-54, 8),
    to_signed(-51, 8),
    to_signed(-38, 8),
    to_signed(-18, 8),
    to_signed(3, 8),
    to_signed(23, 8),
    to_signed(39, 8),
    to_signed(48, 8),
    to_signed(51, 8),
    to_signed(47, 8),
    to_signed(37, 8),
    to_signed(21, 8),
    to_signed(1, 8),
    to_signed(-18, 8),
    to_signed(-33, 8),
    to_signed(-42, 8),
    to_signed(-42, 8),
    to_signed(-34, 8),
    to_signed(-22, 8),
    to_signed(-8, 8),
    to_signed(6, 8),
    to_signed(14, 8),
    to_signed(13, 8),
    to_signed(5, 8),
    to_signed(-8, 8),
    to_signed(-24, 8),
    to_signed(-39, 8),
    to_signed(-51, 8),
    to_signed(-56, 8),
    to_signed(-52, 8),
    to_signed(-38, 8),
    to_signed(-19, 8),
    to_signed(2, 8),
    to_signed(20, 8),
    to_signed(34, 8),
    to_signed(44, 8),
    to_signed(51, 8),
    to_signed(53, 8),
    to_signed(51, 8),
    to_signed(43, 8),
    to_signed(30, 8),
    to_signed(17, 8),
    to_signed(6, 8),
    to_signed(2, 8),
    to_signed(3, 8),
    to_signed(7, 8),
    to_signed(13, 8),
    to_signed(20, 8),
    to_signed(28, 8),
    to_signed(36, 8),
    to_signed(41, 8),
    to_signed(42, 8),
    to_signed(38, 8),
    to_signed(31, 8),
    to_signed(23, 8),
    to_signed(13, 8),
    to_signed(1, 8),
    to_signed(-14, 8),
    to_signed(-34, 8),
    to_signed(-57, 8),
    to_signed(-79, 8),
    to_signed(-91, 8),
    to_signed(-88, 8),
    to_signed(-68, 8),
    to_signed(-37, 8),
    to_signed(-7, 8),
    to_signed(16, 8),
    to_signed(28, 8),
    to_signed(31, 8),
    to_signed(24, 8),
    to_signed(9, 8),
    to_signed(-13, 8),
    to_signed(-36, 8),
    to_signed(-53, 8),
    to_signed(-58, 8),
    to_signed(-50, 8),
    to_signed(-35, 8),
    to_signed(-14, 8),
    to_signed(7, 8),
    to_signed(26, 8),
    to_signed(38, 8),
    to_signed(42, 8),
    to_signed(38, 8),
    to_signed(29, 8),
    to_signed(14, 8),
    to_signed(-3, 8),
    to_signed(-21, 8),
    to_signed(-36, 8),
    to_signed(-43, 8),
    to_signed(-41, 8),
    to_signed(-32, 8),
    to_signed(-19, 8),
    to_signed(-6, 8),
    to_signed(6, 8),
    to_signed(13, 8),
    to_signed(14, 8),
    to_signed(7, 8),
    to_signed(-3, 8),
    to_signed(-16, 8),
    to_signed(-30, 8),
    to_signed(-42, 8),
    to_signed(-49, 8),
    to_signed(-48, 8),
    to_signed(-36, 8),
    to_signed(-17, 8),
    to_signed(6, 8),
    to_signed(26, 8),
    to_signed(40, 8),
    to_signed(50, 8),
    to_signed(57, 8),
    to_signed(60, 8),
    to_signed(59, 8),
    to_signed(53, 8),
    to_signed(40, 8),
    to_signed(25, 8),
    to_signed(10, 8),
    to_signed(0, 8),
    to_signed(-3, 8),
    to_signed(0, 8),
    to_signed(6, 8),
    to_signed(14, 8),
    to_signed(24, 8),
    to_signed(34, 8),
    to_signed(42, 8),
    to_signed(46, 8),
    to_signed(44, 8),
    to_signed(39, 8),
    to_signed(32, 8),
    to_signed(23, 8),
    to_signed(13, 8),
    to_signed(0, 8),
    to_signed(-15, 8),
    to_signed(-33, 8),
    to_signed(-54, 8),
    to_signed(-75, 8),
    to_signed(-87, 8),
    to_signed(-83, 8),
    to_signed(-61, 8),
    to_signed(-30, 8),
    to_signed(-1, 8),
    to_signed(20, 8),
    to_signed(30, 8),
    to_signed(31, 8),
    to_signed(20, 8),
    to_signed(0, 8),
    to_signed(-26, 8),
    to_signed(-50, 8),
    to_signed(-64, 8),
    to_signed(-67, 8),
    to_signed(-59, 8),
    to_signed(-43, 8),
    to_signed(-20, 8),
    to_signed(6, 8),
    to_signed(29, 8),
    to_signed(44, 8),
    to_signed(48, 8),
    to_signed(42, 8),
    to_signed(31, 8),
    to_signed(16, 8),
    to_signed(-3, 8),
    to_signed(-21, 8),
    to_signed(-35, 8),
    to_signed(-41, 8),
    to_signed(-38, 8),
    to_signed(-29, 8),
    to_signed(-18, 8),
    to_signed(-6, 8),
    to_signed(5, 8),
    to_signed(11, 8),
    to_signed(10, 8),
    to_signed(5, 8),
    to_signed(-3, 8),
    to_signed(-12, 8),
    to_signed(-22, 8),
    to_signed(-33, 8),
    to_signed(-40, 8),
    to_signed(-39, 8),
    to_signed(-29, 8),
    to_signed(-12, 8),
    to_signed(9, 8),
    to_signed(28, 8),
    to_signed(44, 8),
    to_signed(56, 8),
    to_signed(61, 8),
    to_signed(61, 8),
    to_signed(56, 8),
    to_signed(47, 8),
    to_signed(36, 8),
    to_signed(23, 8),
    to_signed(11, 8),
    to_signed(2, 8),
    to_signed(0, 8),
    to_signed(2, 8),
    to_signed(6, 8),
    to_signed(12, 8),
    to_signed(22, 8),
    to_signed(33, 8),
    to_signed(44, 8),
    to_signed(51, 8),
    to_signed(52, 8),
    to_signed(50, 8),
    to_signed(44, 8),
    to_signed(34, 8),
    to_signed(19, 8),
    to_signed(0, 8),
    to_signed(-22, 8),
    to_signed(-45, 8),
    to_signed(-68, 8),
    to_signed(-88, 8),
    to_signed(-96, 8),
    to_signed(-89, 8),
    to_signed(-66, 8),
    to_signed(-36, 8),
    to_signed(-7, 8),
    to_signed(15, 8),
    to_signed(29, 8),
    to_signed(35, 8),
    to_signed(28, 8),
    to_signed(9, 8),
    to_signed(-17, 8),
    to_signed(-42, 8),
    to_signed(-58, 8),
    to_signed(-63, 8),
    to_signed(-57, 8),
    to_signed(-42, 8),
    to_signed(-20, 8),
    to_signed(7, 8),
    to_signed(30, 8),
    to_signed(45, 8),
    to_signed(51, 8),
    to_signed(47, 8),
    to_signed(38, 8),
    to_signed(22, 8),
    to_signed(3, 8),
    to_signed(-16, 8),
    to_signed(-28, 8),
    to_signed(-32, 8),
    to_signed(-28, 8),
    to_signed(-21, 8),
    to_signed(-12, 8),
    to_signed(-2, 8),
    to_signed(7, 8),
    to_signed(13, 8),
    to_signed(14, 8),
    to_signed(10, 8),
    to_signed(1, 8),
    to_signed(-11, 8),
    to_signed(-25, 8),
    to_signed(-39, 8),
    to_signed(-49, 8),
    to_signed(-49, 8),
    to_signed(-37, 8),
    to_signed(-17, 8),
    to_signed(6, 8),
    to_signed(28, 8),
    to_signed(45, 8),
    to_signed(55, 8),
    to_signed(59, 8),
    to_signed(59, 8),
    to_signed(53, 8),
    to_signed(43, 8),
    to_signed(30, 8),
    to_signed(16, 8),
    to_signed(5, 8),
    to_signed(-2, 8),
    to_signed(-4, 8),
    to_signed(-3, 8),
    to_signed(0, 8),
    to_signed(7, 8),
    to_signed(17, 8),
    to_signed(28, 8),
    to_signed(37, 8),
    to_signed(43, 8),
    to_signed(44, 8),
    to_signed(42, 8),
    to_signed(36, 8),
    to_signed(25, 8),
    to_signed(10, 8),
    to_signed(-7, 8),
    to_signed(-27, 8),
    to_signed(-47, 8),
    to_signed(-69, 8),
    to_signed(-86, 8),
    to_signed(-94, 8),
    to_signed(-86, 8),
    to_signed(-65, 8),
    to_signed(-36, 8),
    to_signed(-8, 8),
    to_signed(16, 8),
    to_signed(32, 8),
    to_signed(37, 8),
    to_signed(30, 8),
    to_signed(12, 8),
    to_signed(-13, 8),
    to_signed(-37, 8),
    to_signed(-54, 8),
    to_signed(-59, 8),
    to_signed(-54, 8),
    to_signed(-41, 8),
    to_signed(-21, 8),
    to_signed(1, 8),
    to_signed(22, 8),
    to_signed(38, 8),
    to_signed(45, 8),
    to_signed(45, 8),
    to_signed(38, 8),
    to_signed(26, 8),
    to_signed(10, 8),
    to_signed(-5, 8),
    to_signed(-18, 8),
    to_signed(-24, 8),
    to_signed(-25, 8),
    to_signed(-21, 8),
    to_signed(-14, 8),
    to_signed(-7, 8),
    to_signed(0, 8),
    to_signed(4, 8),
    to_signed(5, 8),
    to_signed(3, 8),
    to_signed(-4, 8),
    to_signed(-16, 8),
    to_signed(-31, 8),
    to_signed(-44, 8),
    to_signed(-52, 8),
    to_signed(-51, 8),
    to_signed(-41, 8),
    to_signed(-25, 8),
    to_signed(-5, 8),
    to_signed(15, 8),
    to_signed(32, 8),
    to_signed(44, 8),
    to_signed(52, 8),
    to_signed(54, 8),
    to_signed(50, 8),
    to_signed(42, 8),
    to_signed(29, 8),
    to_signed(15, 8),
    to_signed(4, 8),
    to_signed(-4, 8),
    to_signed(-8, 8),
    to_signed(-8, 8),
    to_signed(-3, 8),
    to_signed(7, 8),
    to_signed(19, 8),
    to_signed(31, 8),
    to_signed(40, 8),
    to_signed(45, 8),
    to_signed(48, 8),
    to_signed(49, 8),
    to_signed(44, 8),
    to_signed(34, 8),
    to_signed(19, 8),
    to_signed(-1, 8),
    to_signed(-23, 8),
    to_signed(-47, 8),
    to_signed(-70, 8),
    to_signed(-87, 8),
    to_signed(-90, 8),
    to_signed(-78, 8),
    to_signed(-52, 8),
    to_signed(-22, 8),
    to_signed(7, 8),
    to_signed(30, 8),
    to_signed(43, 8),
    to_signed(43, 8),
    to_signed(30, 8),
    to_signed(7, 8),
    to_signed(-19, 8),
    to_signed(-39, 8),
    to_signed(-50, 8),
    to_signed(-49, 8),
    to_signed(-39, 8),
    to_signed(-23, 8),
    to_signed(-3, 8),
    to_signed(16, 8),
    to_signed(33, 8),
    to_signed(44, 8),
    to_signed(49, 8),
    to_signed(47, 8),
    to_signed(38, 8),
    to_signed(25, 8),
    to_signed(8, 8),
    to_signed(-9, 8),
    to_signed(-22, 8),
    to_signed(-30, 8),
    to_signed(-30, 8),
    to_signed(-25, 8),
    to_signed(-17, 8),
    to_signed(-10, 8),
    to_signed(-4, 8),
    to_signed(1, 8),
    to_signed(3, 8),
    to_signed(2, 8),
    to_signed(-6, 8),
    to_signed(-20, 8),
    to_signed(-36, 8),
    to_signed(-46, 8),
    to_signed(-47, 8),
    to_signed(-40, 8),
    to_signed(-28, 8),
    to_signed(-12, 8),
    to_signed(6, 8),
    to_signed(25, 8),
    to_signed(41, 8),
    to_signed(53, 8),
    to_signed(58, 8),
    to_signed(57, 8),
    to_signed(52, 8),
    to_signed(42, 8),
    to_signed(28, 8),
    to_signed(14, 8),
    to_signed(2, 8),
    to_signed(-3, 8),
    to_signed(-2, 8),
    to_signed(4, 8),
    to_signed(15, 8),
    to_signed(30, 8),
    to_signed(45, 8),
    to_signed(58, 8),
    to_signed(63, 8),
    to_signed(62, 8),
    to_signed(56, 8),
    to_signed(47, 8),
    to_signed(37, 8),
    to_signed(22, 8),
    to_signed(2, 8),
    to_signed(-21, 8),
    to_signed(-45, 8),
    to_signed(-67, 8),
    to_signed(-83, 8),
    to_signed(-87, 8),
    to_signed(-76, 8),
    to_signed(-51, 8),
    to_signed(-22, 8),
    to_signed(5, 8),
    to_signed(25, 8),
    to_signed(35, 8),
    to_signed(36, 8),
    to_signed(26, 8),
    to_signed(7, 8),
    to_signed(-17, 8),
    to_signed(-39, 8),
    to_signed(-51, 8),
    to_signed(-52, 8),
    to_signed(-43, 8),
    to_signed(-28, 8),
    to_signed(-9, 8),
    to_signed(10, 8),
    to_signed(26, 8),
    to_signed(37, 8),
    to_signed(41, 8),
    to_signed(40, 8),
    to_signed(33, 8),
    to_signed(20, 8),
    to_signed(3, 8),
    to_signed(-15, 8),
    to_signed(-29, 8),
    to_signed(-35, 8),
    to_signed(-33, 8),
    to_signed(-25, 8),
    to_signed(-14, 8),
    to_signed(-3, 8),
    to_signed(6, 8),
    to_signed(11, 8),
    to_signed(10, 8),
    to_signed(5, 8),
    to_signed(-5, 8),
    to_signed(-19, 8),
    to_signed(-34, 8),
    to_signed(-45, 8),
    to_signed(-49, 8),
    to_signed(-44, 8),
    to_signed(-30, 8),
    to_signed(-12, 8),
    to_signed(8, 8),
    to_signed(26, 8),
    to_signed(41, 8),
    to_signed(53, 8),
    to_signed(60, 8),
    to_signed(62, 8),
    to_signed(57, 8),
    to_signed(49, 8),
    to_signed(36, 8),
    to_signed(21, 8),
    to_signed(7, 8),
    to_signed(-2, 8),
    to_signed(-5, 8),
    to_signed(-1, 8),
    to_signed(7, 8),
    to_signed(20, 8),
    to_signed(35, 8),
    to_signed(48, 8),
    to_signed(58, 8),
    to_signed(61, 8),
    to_signed(57, 8),
    to_signed(49, 8),
    to_signed(36, 8),
    to_signed(19, 8),
    to_signed(0, 8),
    to_signed(-23, 8),
    to_signed(-46, 8),
    to_signed(-67, 8),
    to_signed(-84, 8),
    to_signed(-89, 8),
    to_signed(-80, 8),
    to_signed(-58, 8),
    to_signed(-29, 8),
    to_signed(-2, 8),
    to_signed(18, 8),
    to_signed(30, 8),
    to_signed(31, 8),
    to_signed(24, 8),
    to_signed(8, 8),
    to_signed(-14, 8),
    to_signed(-36, 8),
    to_signed(-51, 8),
    to_signed(-56, 8),
    to_signed(-51, 8),
    to_signed(-39, 8),
    to_signed(-21, 8),
    to_signed(0, 8),
    to_signed(22, 8),
    to_signed(38, 8),
    to_signed(46, 8),
    to_signed(46, 8),
    to_signed(40, 8),
    to_signed(28, 8),
    to_signed(12, 8),
    to_signed(-5, 8),
    to_signed(-22, 8),
    to_signed(-34, 8),
    to_signed(-36, 8),
    to_signed(-30, 8),
    to_signed(-19, 8),
    to_signed(-6, 8),
    to_signed(7, 8),
    to_signed(15, 8),
    to_signed(16, 8),
    to_signed(10, 8),
    to_signed(-2, 8),
    to_signed(-17, 8),
    to_signed(-32, 8),
    to_signed(-44, 8),
    to_signed(-49, 8),
    to_signed(-47, 8),
    to_signed(-37, 8),
    to_signed(-19, 8),
    to_signed(4, 8),
    to_signed(24, 8),
    to_signed(39, 8),
    to_signed(48, 8),
    to_signed(54, 8),
    to_signed(57, 8),
    to_signed(55, 8),
    to_signed(47, 8),
    to_signed(33, 8),
    to_signed(17, 8),
    to_signed(3, 8),
    to_signed(-8, 8),
    to_signed(-13, 8),
    to_signed(-14, 8),
    to_signed(-10, 8),
    to_signed(1, 8),
    to_signed(16, 8),
    to_signed(31, 8),
    to_signed(44, 8),
    to_signed(52, 8),
    to_signed(54, 8),
    to_signed(51, 8),
    to_signed(42, 8),
    to_signed(30, 8),
    to_signed(13, 8),
    to_signed(-8, 8),
    to_signed(-31, 8),
    to_signed(-55, 8),
    to_signed(-77, 8),
    to_signed(-91, 8),
    to_signed(-91, 8),
    to_signed(-76, 8),
    to_signed(-50, 8),
    to_signed(-21, 8),
    to_signed(3, 8),
    to_signed(21, 8),
    to_signed(30, 8),
    to_signed(27, 8),
    to_signed(14, 8),
    to_signed(-6, 8),
    to_signed(-29, 8),
    to_signed(-49, 8),
    to_signed(-58, 8),
    to_signed(-58, 8),
    to_signed(-50, 8),
    to_signed(-34, 8),
    to_signed(-13, 8),
    to_signed(8, 8),
    to_signed(26, 8),
    to_signed(37, 8),
    to_signed(42, 8),
    to_signed(40, 8),
    to_signed(32, 8),
    to_signed(19, 8),
    to_signed(5, 8),
    to_signed(-10, 8),
    to_signed(-22, 8),
    to_signed(-29, 8),
    to_signed(-29, 8),
    to_signed(-23, 8),
    to_signed(-13, 8),
    to_signed(-1, 8),
    to_signed(8, 8),
    to_signed(11, 8),
    to_signed(8, 8),
    to_signed(0, 8),
    to_signed(-11, 8),
    to_signed(-23, 8),
    to_signed(-33, 8),
    to_signed(-39, 8),
    to_signed(-40, 8),
    to_signed(-36, 8),
    to_signed(-25, 8),
    to_signed(-10, 8),
    to_signed(8, 8),
    to_signed(23, 8),
    to_signed(34, 8),
    to_signed(42, 8),
    to_signed(47, 8),
    to_signed(48, 8),
    to_signed(46, 8),
    to_signed(40, 8),
    to_signed(30, 8),
    to_signed(18, 8),
    to_signed(9, 8),
    to_signed(2, 8),
    to_signed(-2, 8),
    to_signed(-3, 8),
    to_signed(2, 8),
    to_signed(14, 8),
    to_signed(28, 8),
    to_signed(41, 8),
    to_signed(51, 8),
    to_signed(56, 8),
    to_signed(57, 8),
    to_signed(53, 8),
    to_signed(43, 8),
    to_signed(27, 8),
    to_signed(6, 8),
    to_signed(-19, 8),
    to_signed(-43, 8),
    to_signed(-67, 8),
    to_signed(-85, 8),
    to_signed(-91, 8),
    to_signed(-82, 8),
    to_signed(-58, 8),
    to_signed(-30, 8),
    to_signed(-4, 8),
    to_signed(16, 8),
    to_signed(28, 8),
    to_signed(30, 8),
    to_signed(21, 8),
    to_signed(4, 8),
    to_signed(-19, 8),
    to_signed(-40, 8),
    to_signed(-52, 8),
    to_signed(-53, 8),
    to_signed(-44, 8),
    to_signed(-28, 8),
    to_signed(-7, 8),
    to_signed(16, 8),
    to_signed(34, 8),
    to_signed(46, 8),
    to_signed(49, 8),
    to_signed(44, 8),
    to_signed(32, 8),
    to_signed(16, 8),
    to_signed(0, 8),
    to_signed(-14, 8),
    to_signed(-25, 8),
    to_signed(-32, 8),
    to_signed(-31, 8),
    to_signed(-24, 8),
    to_signed(-12, 8),
    to_signed(1, 8),
    to_signed(12, 8),
    to_signed(17, 8),
    to_signed(13, 8),
    to_signed(3, 8),
    to_signed(-10, 8),
    to_signed(-25, 8),
    to_signed(-39, 8),
    to_signed(-51, 8),
    to_signed(-55, 8),
    to_signed(-52, 8),
    to_signed(-42, 8),
    to_signed(-25, 8),
    to_signed(-6, 8),
    to_signed(13, 8),
    to_signed(29, 8),
    to_signed(42, 8),
    to_signed(50, 8),
    to_signed(53, 8),
    to_signed(51, 8),
    to_signed(45, 8),
    to_signed(35, 8),
    to_signed(23, 8),
    to_signed(12, 8),
    to_signed(5, 8),
    to_signed(3, 8),
    to_signed(4, 8),
    to_signed(9, 8),
    to_signed(18, 8),
    to_signed(32, 8),
    to_signed(45, 8),
    to_signed(54, 8),
    to_signed(57, 8),
    to_signed(53, 8),
    to_signed(44, 8),
    to_signed(33, 8),
    to_signed(18, 8),
    to_signed(0, 8),
    to_signed(-22, 8),
    to_signed(-43, 8),
    to_signed(-63, 8),
    to_signed(-78, 8),
    to_signed(-84, 8),
    to_signed(-77, 8),
    to_signed(-57, 8),
    to_signed(-30, 8),
    to_signed(-4, 8),
    to_signed(16, 8),
    to_signed(28, 8),
    to_signed(28, 8),
    to_signed(19, 8),
    to_signed(0, 8),
    to_signed(-23, 8),
    to_signed(-45, 8),
    to_signed(-57, 8),
    to_signed(-57, 8),
    to_signed(-48, 8),
    to_signed(-32, 8),
    to_signed(-12, 8),
    to_signed(10, 8),
    to_signed(30, 8),
    to_signed(43, 8),
    to_signed(46, 8),
    to_signed(40, 8),
    to_signed(28, 8),
    to_signed(12, 8),
    to_signed(-4, 8),
    to_signed(-18, 8),
    to_signed(-29, 8),
    to_signed(-36, 8),
    to_signed(-37, 8),
    to_signed(-31, 8),
    to_signed(-19, 8),
    to_signed(-5, 8),
    to_signed(6, 8),
    to_signed(10, 8),
    to_signed(6, 8),
    to_signed(-3, 8),
    to_signed(-13, 8),
    to_signed(-25, 8),
    to_signed(-39, 8),
    to_signed(-50, 8),
    to_signed(-54, 8),
    to_signed(-49, 8),
    to_signed(-37, 8),
    to_signed(-19, 8),
    to_signed(0, 8),
    to_signed(20, 8),
    to_signed(36, 8),
    to_signed(47, 8),
    to_signed(55, 8),
    to_signed(57, 8),
    to_signed(54, 8),
    to_signed(49, 8),
    to_signed(40, 8),
    to_signed(28, 8),
    to_signed(16, 8),
    to_signed(9, 8),
    to_signed(7, 8),
    to_signed(8, 8),
    to_signed(11, 8),
    to_signed(17, 8),
    to_signed(26, 8),
    to_signed(36, 8),
    to_signed(44, 8),
    to_signed(47, 8),
    to_signed(46, 8),
    to_signed(40, 8),
    to_signed(33, 8),
    to_signed(23, 8),
    to_signed(10, 8),
    to_signed(-9, 8),
    to_signed(-31, 8),
    to_signed(-53, 8),
    to_signed(-71, 8),
    to_signed(-81, 8),
    to_signed(-79, 8),
    to_signed(-64, 8),
    to_signed(-39, 8),
    to_signed(-13, 8),
    to_signed(11, 8),
    to_signed(28, 8),
    to_signed(34, 8),
    to_signed(28, 8),
    to_signed(9, 8),
    to_signed(-15, 8),
    to_signed(-38, 8),
    to_signed(-54, 8),
    to_signed(-59, 8),
    to_signed(-54, 8),
    to_signed(-43, 8),
    to_signed(-26, 8),
    to_signed(-4, 8),
    to_signed(18, 8),
    to_signed(35, 8),
    to_signed(44, 8),
    to_signed(46, 8),
    to_signed(40, 8),
    to_signed(28, 8),
    to_signed(11, 8),
    to_signed(-7, 8),
    to_signed(-24, 8),
    to_signed(-36, 8),
    to_signed(-42, 8),
    to_signed(-39, 8),
    to_signed(-31, 8),
    to_signed(-19, 8),
    to_signed(-7, 8),
    to_signed(2, 8),
    to_signed(7, 8),
    to_signed(5, 8),
    to_signed(-1, 8),
    to_signed(-10, 8),
    to_signed(-21, 8),
    to_signed(-33, 8),
    to_signed(-40, 8),
    to_signed(-41, 8),
    to_signed(-35, 8),
    to_signed(-24, 8),
    to_signed(-10, 8),
    to_signed(5, 8),
    to_signed(19, 8),
    to_signed(30, 8),
    to_signed(40, 8),
    to_signed(46, 8),
    to_signed(48, 8),
    to_signed(45, 8),
    to_signed(38, 8),
    to_signed(29, 8),
    to_signed(19, 8),
    to_signed(11, 8),
    to_signed(7, 8),
    to_signed(6, 8),
    to_signed(7, 8),
    to_signed(12, 8),
    to_signed(23, 8),
    to_signed(35, 8),
    to_signed(47, 8),
    to_signed(54, 8),
    to_signed(58, 8),
    to_signed(58, 8),
    to_signed(54, 8),
    to_signed(44, 8),
    to_signed(29, 8),
    to_signed(7, 8),
    to_signed(-19, 8),
    to_signed(-46, 8),
    to_signed(-70, 8),
    to_signed(-88, 8),
    to_signed(-92, 8),
    to_signed(-79, 8),
    to_signed(-52, 8),
    to_signed(-21, 8),
    to_signed(5, 8),
    to_signed(24, 8),
    to_signed(31, 8),
    to_signed(28, 8),
    to_signed(14, 8),
    to_signed(-9, 8),
    to_signed(-35, 8),
    to_signed(-55, 8),
    to_signed(-64, 8),
    to_signed(-59, 8),
    to_signed(-48, 8),
    to_signed(-31, 8),
    to_signed(-11, 8),
    to_signed(10, 8),
    to_signed(28, 8),
    to_signed(39, 8),
    to_signed(41, 8),
    to_signed(37, 8),
    to_signed(28, 8),
    to_signed(16, 8),
    to_signed(1, 8),
    to_signed(-16, 8),
    to_signed(-32, 8),
    to_signed(-41, 8),
    to_signed(-40, 8),
    to_signed(-31, 8),
    to_signed(-18, 8),
    to_signed(-5, 8),
    to_signed(4, 8),
    to_signed(9, 8),
    to_signed(8, 8),
    to_signed(1, 8),
    to_signed(-10, 8),
    to_signed(-23, 8),
    to_signed(-34, 8),
    to_signed(-40, 8),
    to_signed(-38, 8),
    to_signed(-33, 8),
    to_signed(-24, 8),
    to_signed(-11, 8),
    to_signed(5, 8),
    to_signed(21, 8),
    to_signed(35, 8),
    to_signed(45, 8),
    to_signed(52, 8),
    to_signed(56, 8),
    to_signed(57, 8),
    to_signed(53, 8),
    to_signed(45, 8),
    to_signed(33, 8),
    to_signed(22, 8),
    to_signed(16, 8),
    to_signed(15, 8),
    to_signed(17, 8),
    to_signed(23, 8),
    to_signed(30, 8),
    to_signed(40, 8),
    to_signed(47, 8),
    to_signed(53, 8),
    to_signed(54, 8),
    to_signed(52, 8),
    to_signed(45, 8),
    to_signed(34, 8),
    to_signed(19, 8),
    to_signed(-2, 8),
    to_signed(-27, 8),
    to_signed(-52, 8),
    to_signed(-73, 8),
    to_signed(-87, 8),
    to_signed(-87, 8),
    to_signed(-72, 8),
    to_signed(-46, 8),
    to_signed(-17, 8),
    to_signed(8, 8),
    to_signed(25, 8),
    to_signed(30, 8),
    to_signed(24, 8),
    to_signed(9, 8),
    to_signed(-13, 8),
    to_signed(-34, 8),
    to_signed(-51, 8),
    to_signed(-57, 8),
    to_signed(-52, 8),
    to_signed(-39, 8),
    to_signed(-23, 8),
    to_signed(-5, 8),
    to_signed(13, 8),
    to_signed(28, 8),
    to_signed(38, 8),
    to_signed(41, 8),
    to_signed(38, 8),
    to_signed(28, 8),
    to_signed(14, 8),
    to_signed(-2, 8),
    to_signed(-17, 8),
    to_signed(-31, 8),
    to_signed(-40, 8),
    to_signed(-41, 8),
    to_signed(-32, 8),
    to_signed(-19, 8),
    to_signed(-6, 8),
    to_signed(3, 8),
    to_signed(6, 8),
    to_signed(3, 8),
    to_signed(-5, 8),
    to_signed(-16, 8),
    to_signed(-27, 8),
    to_signed(-36, 8),
    to_signed(-39, 8),
    to_signed(-36, 8),
    to_signed(-28, 8),
    to_signed(-19, 8),
    to_signed(-8, 8),
    to_signed(6, 8),
    to_signed(21, 8),
    to_signed(35, 8),
    to_signed(47, 8),
    to_signed(54, 8),
    to_signed(59, 8),
    to_signed(58, 8),
    to_signed(53, 8),
    to_signed(43, 8),
    to_signed(30, 8),
    to_signed(17, 8),
    to_signed(8, 8),
    to_signed(6, 8),
    to_signed(9, 8),
    to_signed(17, 8),
    to_signed(27, 8),
    to_signed(38, 8),
    to_signed(46, 8),
    to_signed(50, 8),
    to_signed(48, 8),
    to_signed(42, 8),
    to_signed(32, 8),
    to_signed(19, 8),
    to_signed(3, 8),
    to_signed(-16, 8),
    to_signed(-39, 8),
    to_signed(-61, 8),
    to_signed(-79, 8),
    to_signed(-86, 8),
    to_signed(-81, 8),
    to_signed(-62, 8),
    to_signed(-36, 8),
    to_signed(-11, 8),
    to_signed(10, 8),
    to_signed(22, 8),
    to_signed(23, 8),
    to_signed(14, 8),
    to_signed(-4, 8),
    to_signed(-27, 8),
    to_signed(-47, 8),
    to_signed(-59, 8),
    to_signed(-60, 8),
    to_signed(-50, 8),
    to_signed(-33, 8),
    to_signed(-13, 8),
    to_signed(7, 8),
    to_signed(25, 8),
    to_signed(39, 8),
    to_signed(47, 8),
    to_signed(48, 8),
    to_signed(42, 8),
    to_signed(29, 8),
    to_signed(13, 8),
    to_signed(-6, 8),
    to_signed(-22, 8),
    to_signed(-35, 8),
    to_signed(-40, 8),
    to_signed(-36, 8),
    to_signed(-24, 8),
    to_signed(-8, 8),
    to_signed(5, 8),
    to_signed(13, 8),
    to_signed(13, 8),
    to_signed(6, 8),
    to_signed(-5, 8),
    to_signed(-17, 8),
    to_signed(-28, 8),
    to_signed(-34, 8),
    to_signed(-34, 8),
    to_signed(-27, 8),
    to_signed(-15, 8),
    to_signed(-1, 8),
    to_signed(12, 8),
    to_signed(25, 8),
    to_signed(36, 8),
    to_signed(46, 8),
    to_signed(52, 8),
    to_signed(55, 8),
    to_signed(54, 8),
    to_signed(49, 8),
    to_signed(40, 8),
    to_signed(29, 8),
    to_signed(16, 8),
    to_signed(7, 8),
    to_signed(3, 8),
    to_signed(6, 8),
    to_signed(15, 8),
    to_signed(27, 8),
    to_signed(41, 8),
    to_signed(53, 8),
    to_signed(61, 8),
    to_signed(60, 8),
    to_signed(52, 8),
    to_signed(38, 8),
    to_signed(21, 8),
    to_signed(3, 8),
    to_signed(-16, 8),
    to_signed(-37, 8),
    to_signed(-59, 8),
    to_signed(-76, 8),
    to_signed(-85, 8),
    to_signed(-81, 8),
    to_signed(-67, 8),
    to_signed(-44, 8),
    to_signed(-18, 8),
    to_signed(5, 8),
    to_signed(20, 8),
    to_signed(25, 8),
    to_signed(19, 8),
    to_signed(3, 8),
    to_signed(-19, 8),
    to_signed(-41, 8),
    to_signed(-56, 8),
    to_signed(-59, 8),
    to_signed(-51, 8),
    to_signed(-35, 8),
    to_signed(-14, 8),
    to_signed(7, 8),
    to_signed(25, 8),
    to_signed(39, 8),
    to_signed(47, 8),
    to_signed(49, 8),
    to_signed(43, 8),
    to_signed(33, 8),
    to_signed(19, 8),
    to_signed(4, 8),
    to_signed(-12, 8),
    to_signed(-27, 8),
    to_signed(-35, 8),
    to_signed(-35, 8),
    to_signed(-26, 8),
    to_signed(-9, 8),
    to_signed(8, 8),
    to_signed(21, 8),
    to_signed(26, 8),
    to_signed(22, 8),
    to_signed(9, 8),
    to_signed(-9, 8),
    to_signed(-28, 8),
    to_signed(-42, 8),
    to_signed(-48, 8),
    to_signed(-44, 8),
    to_signed(-33, 8),
    to_signed(-16, 8),
    to_signed(2, 8),
    to_signed(18, 8),
    to_signed(29, 8),
    to_signed(36, 8),
    to_signed(40, 8),
    to_signed(43, 8),
    to_signed(43, 8),
    to_signed(39, 8),
    to_signed(32, 8),
    to_signed(22, 8),
    to_signed(13, 8),
    to_signed(5, 8),
    to_signed(-1, 8),
    to_signed(-2, 8),
    to_signed(3, 8),
    to_signed(14, 8),
    to_signed(30, 8),
    to_signed(45, 8),
    to_signed(55, 8),
    to_signed(59, 8),
    to_signed(55, 8),
    to_signed(44, 8),
    to_signed(25, 8),
    to_signed(3, 8),
    to_signed(-20, 8),
    to_signed(-42, 8),
    to_signed(-62, 8),
    to_signed(-79, 8),
    to_signed(-90, 8),
    to_signed(-89, 8),
    to_signed(-75, 8),
    to_signed(-52, 8),
    to_signed(-25, 8),
    to_signed(0, 8),
    to_signed(19, 8),
    to_signed(29, 8),
    to_signed(26, 8),
    to_signed(11, 8),
    to_signed(-13, 8),
    to_signed(-36, 8),
    to_signed(-53, 8),
    to_signed(-60, 8),
    to_signed(-56, 8),
    to_signed(-41, 8),
    to_signed(-20, 8),
    to_signed(3, 8),
    to_signed(24, 8),
    to_signed(39, 8),
    to_signed(47, 8),
    to_signed(48, 8),
    to_signed(43, 8),
    to_signed(32, 8),
    to_signed(18, 8),
    to_signed(4, 8),
    to_signed(-8, 8),
    to_signed(-19, 8),
    to_signed(-28, 8),
    to_signed(-31, 8),
    to_signed(-26, 8),
    to_signed(-11, 8),
    to_signed(6, 8),
    to_signed(19, 8),
    to_signed(25, 8),
    to_signed(22, 8),
    to_signed(11, 8),
    to_signed(-6, 8),
    to_signed(-28, 8),
    to_signed(-47, 8),
    to_signed(-58, 8),
    to_signed(-55, 8),
    to_signed(-42, 8),
    to_signed(-21, 8),
    to_signed(1, 8),
    to_signed(22, 8),
    to_signed(38, 8),
    to_signed(46, 8),
    to_signed(48, 8),
    to_signed(45, 8),
    to_signed(41, 8),
    to_signed(38, 8),
    to_signed(32, 8),
    to_signed(24, 8),
    to_signed(15, 8),
    to_signed(8, 8),
    to_signed(3, 8),
    to_signed(2, 8),
    to_signed(4, 8),
    to_signed(11, 8),
    to_signed(24, 8),
    to_signed(39, 8),
    to_signed(51, 8),
    to_signed(56, 8),
    to_signed(53, 8),
    to_signed(44, 8),
    to_signed(29, 8),
    to_signed(10, 8),
    to_signed(-12, 8),
    to_signed(-32, 8),
    to_signed(-50, 8),
    to_signed(-65, 8),
    to_signed(-78, 8),
    to_signed(-84, 8),
    to_signed(-80, 8),
    to_signed(-63, 8),
    to_signed(-40, 8),
    to_signed(-16, 8),
    to_signed(3, 8),
    to_signed(17, 8),
    to_signed(22, 8),
    to_signed(16, 8),
    to_signed(-1, 8),
    to_signed(-26, 8),
    to_signed(-48, 8),
    to_signed(-60, 8),
    to_signed(-59, 8),
    to_signed(-50, 8),
    to_signed(-33, 8),
    to_signed(-12, 8),
    to_signed(10, 8),
    to_signed(30, 8),
    to_signed(42, 8),
    to_signed(45, 8),
    to_signed(41, 8),
    to_signed(35, 8),
    to_signed(25, 8),
    to_signed(12, 8),
    to_signed(-3, 8),
    to_signed(-17, 8),
    to_signed(-28, 8),
    to_signed(-35, 8),
    to_signed(-37, 8),
    to_signed(-32, 8),
    to_signed(-20, 8),
    to_signed(-6, 8),
    to_signed(4, 8),
    to_signed(8, 8),
    to_signed(3, 8),
    to_signed(-8, 8),
    to_signed(-24, 8),
    to_signed(-42, 8),
    to_signed(-57, 8),
    to_signed(-62, 8),
    to_signed(-55, 8),
    to_signed(-38, 8),
    to_signed(-17, 8),
    to_signed(4, 8),
    to_signed(23, 8),
    to_signed(36, 8),
    to_signed(41, 8),
    to_signed(38, 8),
    to_signed(31, 8),
    to_signed(25, 8),
    to_signed(22, 8),
    to_signed(18, 8),
    to_signed(12, 8),
    to_signed(5, 8),
    to_signed(0, 8),
    to_signed(-2, 8),
    to_signed(-1, 8),
    to_signed(1, 8),
    to_signed(5, 8),
    to_signed(15, 8),
    to_signed(29, 8),
    to_signed(42, 8),
    to_signed(48, 8),
    to_signed(47, 8),
    to_signed(41, 8),
    to_signed(32, 8),
    to_signed(18, 8),
    to_signed(1, 8),
    to_signed(-18, 8),
    to_signed(-36, 8),
    to_signed(-53, 8),
    to_signed(-67, 8),
    to_signed(-77, 8),
    to_signed(-77, 8),
    to_signed(-62, 8),
    to_signed(-38, 8),
    to_signed(-11, 8),
    to_signed(10, 8),
    to_signed(25, 8),
    to_signed(32, 8),
    to_signed(29, 8),
    to_signed(15, 8),
    to_signed(-8, 8),
    to_signed(-32, 8),
    to_signed(-47, 8),
    to_signed(-52, 8),
    to_signed(-46, 8),
    to_signed(-34, 8),
    to_signed(-17, 8),
    to_signed(4, 8),
    to_signed(23, 8),
    to_signed(37, 8),
    to_signed(43, 8),
    to_signed(43, 8),
    to_signed(40, 8),
    to_signed(33, 8),
    to_signed(22, 8),
    to_signed(7, 8),
    to_signed(-10, 8),
    to_signed(-24, 8),
    to_signed(-34, 8),
    to_signed(-37, 8),
    to_signed(-34, 8),
    to_signed(-22, 8),
    to_signed(-7, 8),
    to_signed(8, 8),
    to_signed(16, 8),
    to_signed(15, 8),
    to_signed(7, 8),
    to_signed(-7, 8),
    to_signed(-24, 8),
    to_signed(-38, 8),
    to_signed(-47, 8),
    to_signed(-45, 8),
    to_signed(-34, 8),
    to_signed(-18, 8),
    to_signed(0, 8),
    to_signed(18, 8),
    to_signed(33, 8),
    to_signed(42, 8),
    to_signed(44, 8),
    to_signed(42, 8),
    to_signed(39, 8),
    to_signed(37, 8),
    to_signed(34, 8),
    to_signed(29, 8),
    to_signed(21, 8),
    to_signed(14, 8),
    to_signed(10, 8),
    to_signed(9, 8),
    to_signed(12, 8),
    to_signed(17, 8),
    to_signed(29, 8),
    to_signed(44, 8),
    to_signed(58, 8),
    to_signed(67, 8),
    to_signed(67, 8),
    to_signed(61, 8),
    to_signed(50, 8),
    to_signed(34, 8),
    to_signed(14, 8),
    to_signed(-10, 8),
    to_signed(-34, 8),
    to_signed(-56, 8),
    to_signed(-74, 8),
    to_signed(-83, 8),
    to_signed(-78, 8),
    to_signed(-57, 8),
    to_signed(-27, 8),
    to_signed(4, 8),
    to_signed(27, 8),
    to_signed(41, 8),
    to_signed(45, 8),
    to_signed(38, 8),
    to_signed(20, 8),
    to_signed(-8, 8),
    to_signed(-36, 8),
    to_signed(-53, 8),
    to_signed(-56, 8),
    to_signed(-46, 8),
    to_signed(-31, 8),
    to_signed(-12, 8),
    to_signed(9, 8),
    to_signed(29, 8),
    to_signed(44, 8),
    to_signed(51, 8),
    to_signed(50, 8),
    to_signed(43, 8),
    to_signed(33, 8),
    to_signed(19, 8),
    to_signed(3, 8),
    to_signed(-13, 8),
    to_signed(-27, 8),
    to_signed(-36, 8),
    to_signed(-37, 8),
    to_signed(-30, 8),
    to_signed(-17, 8),
    to_signed(0, 8),
    to_signed(14, 8),
    to_signed(20, 8),
    to_signed(17, 8),
    to_signed(4, 8),
    to_signed(-14, 8),
    to_signed(-34, 8),
    to_signed(-50, 8),
    to_signed(-58, 8),
    to_signed(-55, 8),
    to_signed(-43, 8),
    to_signed(-25, 8),
    to_signed(-4, 8),
    to_signed(18, 8),
    to_signed(36, 8),
    to_signed(47, 8),
    to_signed(51, 8),
    to_signed(50, 8),
    to_signed(47, 8),
    to_signed(44, 8),
    to_signed(39, 8),
    to_signed(31, 8),
    to_signed(22, 8),
    to_signed(15, 8),
    to_signed(12, 8),
    to_signed(12, 8),
    to_signed(15, 8),
    to_signed(22, 8),
    to_signed(34, 8),
    to_signed(51, 8),
    to_signed(65, 8),
    to_signed(72, 8),
    to_signed(69, 8),
    to_signed(57, 8),
    to_signed(42, 8),
    to_signed(22, 8),
    to_signed(0, 8),
    to_signed(-24, 8),
    to_signed(-50, 8),
    to_signed(-72, 8),
    to_signed(-86, 8),
    to_signed(-86, 8),
    to_signed(-72, 8),
    to_signed(-45, 8),
    to_signed(-14, 8),
    to_signed(12, 8),
    to_signed(29, 8),
    to_signed(36, 8),
    to_signed(33, 8),
    to_signed(18, 8),
    to_signed(-9, 8),
    to_signed(-40, 8),
    to_signed(-64, 8),
    to_signed(-73, 8),
    to_signed(-67, 8),
    to_signed(-51, 8),
    to_signed(-30, 8),
    to_signed(-8, 8),
    to_signed(14, 8),
    to_signed(32, 8),
    to_signed(45, 8),
    to_signed(49, 8),
    to_signed(45, 8),
    to_signed(34, 8),
    to_signed(20, 8),
    to_signed(5, 8),
    to_signed(-10, 8),
    to_signed(-24, 8),
    to_signed(-34, 8),
    to_signed(-40, 8),
    to_signed(-39, 8),
    to_signed(-30, 8),
    to_signed(-16, 8),
    to_signed(0, 8),
    to_signed(9, 8),
    to_signed(9, 8),
    to_signed(0, 8),
    to_signed(-14, 8),
    to_signed(-30, 8),
    to_signed(-46, 8),
    to_signed(-57, 8),
    to_signed(-59, 8),
    to_signed(-50, 8),
    to_signed(-33, 8),
    to_signed(-11, 8),
    to_signed(10, 8),
    to_signed(29, 8),
    to_signed(42, 8),
    to_signed(48, 8),
    to_signed(48, 8),
    to_signed(44, 8),
    to_signed(39, 8),
    to_signed(33, 8),
    to_signed(25, 8),
    to_signed(16, 8),
    to_signed(8, 8),
    to_signed(3, 8),
    to_signed(4, 8),
    to_signed(7, 8),
    to_signed(13, 8),
    to_signed(24, 8),
    to_signed(39, 8),
    to_signed(55, 8),
    to_signed(66, 8),
    to_signed(68, 8),
    to_signed(62, 8),
    to_signed(50, 8),
    to_signed(33, 8),
    to_signed(12, 8),
    to_signed(-11, 8),
    to_signed(-34, 8),
    to_signed(-56, 8),
    to_signed(-75, 8),
    to_signed(-87, 8),
    to_signed(-88, 8),
    to_signed(-73, 8),
    to_signed(-47, 8),
    to_signed(-19, 8),
    to_signed(4, 8),
    to_signed(18, 8),
    to_signed(24, 8),
    to_signed(21, 8),
    to_signed(7, 8),
    to_signed(-18, 8),
    to_signed(-48, 8),
    to_signed(-69, 8),
    to_signed(-73, 8),
    to_signed(-61, 8),
    to_signed(-42, 8),
    to_signed(-23, 8),
    to_signed(-4, 8),
    to_signed(16, 8),
    to_signed(32, 8),
    to_signed(42, 8),
    to_signed(41, 8),
    to_signed(32, 8),
    to_signed(21, 8),
    to_signed(8, 8),
    to_signed(-5, 8),
    to_signed(-18, 8),
    to_signed(-30, 8),
    to_signed(-38, 8),
    to_signed(-41, 8),
    to_signed(-37, 8),
    to_signed(-27, 8),
    to_signed(-12, 8),
    to_signed(1, 8),
    to_signed(7, 8),
    to_signed(4, 8),
    to_signed(-5, 8),
    to_signed(-18, 8),
    to_signed(-31, 8),
    to_signed(-43, 8),
    to_signed(-51, 8),
    to_signed(-50, 8),
    to_signed(-39, 8),
    to_signed(-20, 8),
    to_signed(-1, 8),
    to_signed(15, 8),
    to_signed(27, 8),
    to_signed(34, 8),
    to_signed(38, 8),
    to_signed(38, 8),
    to_signed(36, 8),
    to_signed(33, 8),
    to_signed(30, 8),
    to_signed(27, 8),
    to_signed(21, 8),
    to_signed(15, 8),
    to_signed(11, 8),
    to_signed(10, 8),
    to_signed(12, 8),
    to_signed(16, 8),
    to_signed(24, 8),
    to_signed(37, 8),
    to_signed(51, 8),
    to_signed(60, 8),
    to_signed(63, 8),
    to_signed(59, 8),
    to_signed(51, 8),
    to_signed(39, 8),
    to_signed(21, 8),
    to_signed(-1, 8),
    to_signed(-26, 8),
    to_signed(-50, 8),
    to_signed(-70, 8),
    to_signed(-84, 8),
    to_signed(-87, 8),
    to_signed(-76, 8),
    to_signed(-52, 8),
    to_signed(-21, 8),
    to_signed(8, 8),
    to_signed(28, 8),
    to_signed(39, 8),
    to_signed(40, 8),
    to_signed(30, 8),
    to_signed(7, 8),
    to_signed(-22, 8),
    to_signed(-47, 8),
    to_signed(-59, 8),
    to_signed(-56, 8),
    to_signed(-45, 8),
    to_signed(-29, 8),
    to_signed(-10, 8),
    to_signed(11, 8),
    to_signed(32, 8),
    to_signed(47, 8),
    to_signed(52, 8),
    to_signed(50, 8),
    to_signed(44, 8),
    to_signed(36, 8),
    to_signed(24, 8),
    to_signed(9, 8),
    to_signed(-8, 8),
    to_signed(-21, 8),
    to_signed(-27, 8),
    to_signed(-24, 8),
    to_signed(-14, 8),
    to_signed(-2, 8),
    to_signed(11, 8),
    to_signed(18, 8),
    to_signed(19, 8),
    to_signed(11, 8),
    to_signed(-2, 8),
    to_signed(-18, 8),
    to_signed(-33, 8),
    to_signed(-43, 8),
    to_signed(-43, 8),
    to_signed(-34, 8),
    to_signed(-18, 8),
    to_signed(-1, 8),
    to_signed(13, 8),
    to_signed(24, 8),
    to_signed(33, 8),
    to_signed(40, 8),
    to_signed(44, 8),
    to_signed(45, 8),
    to_signed(44, 8),
    to_signed(42, 8),
    to_signed(38, 8),
    to_signed(33, 8),
    to_signed(25, 8),
    to_signed(17, 8),
    to_signed(9, 8),
    to_signed(5, 8),
    to_signed(7, 8),
    to_signed(14, 8),
    to_signed(25, 8),
    to_signed(38, 8),
    to_signed(48, 8),
    to_signed(54, 8),
    to_signed(55, 8),
    to_signed(52, 8),
    to_signed(43, 8),
    to_signed(27, 8),
    to_signed(6, 8),
    to_signed(-18, 8),
    to_signed(-44, 8),
    to_signed(-68, 8),
    to_signed(-87, 8),
    to_signed(-96, 8),
    to_signed(-89, 8),
    to_signed(-67, 8),
    to_signed(-36, 8),
    to_signed(-5, 8),
    to_signed(18, 8),
    to_signed(31, 8),
    to_signed(33, 8),
    to_signed(25, 8),
    to_signed(5, 8),
    to_signed(-21, 8),
    to_signed(-47, 8),
    to_signed(-65, 8),
    to_signed(-70, 8),
    to_signed(-62, 8),
    to_signed(-47, 8),
    to_signed(-26, 8),
    to_signed(-2, 8),
    to_signed(20, 8),
    to_signed(38, 8),
    to_signed(48, 8),
    to_signed(50, 8),
    to_signed(46, 8),
    to_signed(38, 8),
    to_signed(24, 8),
    to_signed(6, 8),
    to_signed(-14, 8),
    to_signed(-30, 8),
    to_signed(-39, 8),
    to_signed(-38, 8),
    to_signed(-29, 8),
    to_signed(-16, 8),
    to_signed(-3, 8),
    to_signed(7, 8),
    to_signed(12, 8),
    to_signed(9, 8),
    to_signed(-1, 8),
    to_signed(-16, 8),
    to_signed(-31, 8),
    to_signed(-41, 8),
    to_signed(-42, 8),
    to_signed(-35, 8),
    to_signed(-23, 8),
    to_signed(-9, 8),
    to_signed(4, 8),
    to_signed(18, 8),
    to_signed(30, 8),
    to_signed(39, 8),
    to_signed(44, 8),
    to_signed(45, 8),
    to_signed(46, 8),
    to_signed(44, 8),
    to_signed(40, 8),
    to_signed(32, 8),
    to_signed(20, 8),
    to_signed(7, 8),
    to_signed(-2, 8),
    to_signed(-4, 8),
    to_signed(0, 8),
    to_signed(11, 8),
    to_signed(26, 8),
    to_signed(42, 8),
    to_signed(57, 8),
    to_signed(66, 8),
    to_signed(68, 8),
    to_signed(62, 8),
    to_signed(49, 8),
    to_signed(29, 8),
    to_signed(5, 8),
    to_signed(-21, 8),
    to_signed(-48, 8),
    to_signed(-73, 8),
    to_signed(-92, 8),
    to_signed(-100, 8),
    to_signed(-92, 8),
    to_signed(-69, 8),
    to_signed(-37, 8),
    to_signed(-6, 8),
    to_signed(18, 8),
    to_signed(31, 8),
    to_signed(34, 8),
    to_signed(26, 8),
    to_signed(6, 8),
    to_signed(-20, 8),
    to_signed(-47, 8),
    to_signed(-66, 8),
    to_signed(-72, 8),
    to_signed(-65, 8),
    to_signed(-47, 8),
    to_signed(-24, 8),
    to_signed(2, 8),
    to_signed(25, 8),
    to_signed(41, 8),
    to_signed(50, 8),
    to_signed(51, 8),
    to_signed(43, 8),
    to_signed(28, 8),
    to_signed(9, 8),
    to_signed(-13, 8),
    to_signed(-30, 8),
    to_signed(-42, 8),
    to_signed(-45, 8),
    to_signed(-40, 8),
    to_signed(-27, 8),
    to_signed(-9, 8),
    to_signed(7, 8),
    to_signed(18, 8),
    to_signed(19, 8),
    to_signed(10, 8),
    to_signed(-5, 8),
    to_signed(-23, 8),
    to_signed(-40, 8),
    to_signed(-51, 8),
    to_signed(-54, 8),
    to_signed(-47, 8),
    to_signed(-33, 8),
    to_signed(-15, 8),
    to_signed(4, 8),
    to_signed(21, 8),
    to_signed(35, 8),
    to_signed(44, 8),
    to_signed(47, 8),
    to_signed(46, 8),
    to_signed(43, 8),
    to_signed(39, 8),
    to_signed(34, 8),
    to_signed(27, 8),
    to_signed(16, 8),
    to_signed(7, 8),
    to_signed(2, 8),
    to_signed(4, 8),
    to_signed(12, 8),
    to_signed(24, 8),
    to_signed(39, 8),
    to_signed(52, 8),
    to_signed(63, 8),
    to_signed(68, 8),
    to_signed(66, 8),
    to_signed(57, 8),
    to_signed(43, 8),
    to_signed(23, 8),
    to_signed(0, 8),
    to_signed(-24, 8),
    to_signed(-47, 8),
    to_signed(-69, 8),
    to_signed(-86, 8),
    to_signed(-93, 8),
    to_signed(-87, 8),
    to_signed(-66, 8),
    to_signed(-38, 8),
    to_signed(-9, 8),
    to_signed(14, 8),
    to_signed(29, 8),
    to_signed(36, 8),
    to_signed(32, 8),
    to_signed(16, 8),
    to_signed(-11, 8),
    to_signed(-41, 8),
    to_signed(-63, 8),
    to_signed(-71, 8),
    to_signed(-66, 8),
    to_signed(-51, 8),
    to_signed(-31, 8),
    to_signed(-8, 8),
    to_signed(15, 8),
    to_signed(35, 8),
    to_signed(48, 8),
    to_signed(52, 8),
    to_signed(47, 8),
    to_signed(35, 8),
    to_signed(17, 8),
    to_signed(-2, 8),
    to_signed(-21, 8),
    to_signed(-34, 8),
    to_signed(-40, 8),
    to_signed(-38, 8),
    to_signed(-28, 8),
    to_signed(-14, 8),
    to_signed(1, 8),
    to_signed(12, 8),
    to_signed(16, 8),
    to_signed(11, 8),
    to_signed(-1, 8),
    to_signed(-16, 8),
    to_signed(-33, 8),
    to_signed(-46, 8),
    to_signed(-53, 8),
    to_signed(-52, 8),
    to_signed(-41, 8),
    to_signed(-25, 8),
    to_signed(-6, 8),
    to_signed(13, 8),
    to_signed(29, 8),
    to_signed(40, 8),
    to_signed(48, 8),
    to_signed(50, 8),
    to_signed(50, 8),
    to_signed(46, 8),
    to_signed(40, 8),
    to_signed(32, 8),
    to_signed(21, 8),
    to_signed(11, 8),
    to_signed(6, 8),
    to_signed(7, 8),
    to_signed(13, 8),
    to_signed(21, 8),
    to_signed(32, 8),
    to_signed(43, 8),
    to_signed(54, 8),
    to_signed(63, 8),
    to_signed(66, 8),
    to_signed(63, 8),
    to_signed(53, 8),
    to_signed(38, 8),
    to_signed(19, 8),
    to_signed(-4, 8),
    to_signed(-30, 8),
    to_signed(-56, 8),
    to_signed(-78, 8),
    to_signed(-92, 8),
    to_signed(-91, 8),
    to_signed(-76, 8),
    to_signed(-49, 8),
    to_signed(-18, 8),
    to_signed(10, 8),
    to_signed(30, 8),
    to_signed(40, 8),
    to_signed(36, 8),
    to_signed(20, 8),
    to_signed(-7, 8),
    to_signed(-37, 8),
    to_signed(-62, 8),
    to_signed(-75, 8),
    to_signed(-74, 8),
    to_signed(-61, 8),
    to_signed(-39, 8),
    to_signed(-13, 8),
    to_signed(13, 8),
    to_signed(35, 8),
    to_signed(49, 8),
    to_signed(54, 8),
    to_signed(51, 8),
    to_signed(42, 8),
    to_signed(27, 8),
    to_signed(10, 8),
    to_signed(-9, 8),
    to_signed(-26, 8),
    to_signed(-38, 8),
    to_signed(-40, 8),
    to_signed(-34, 8),
    to_signed(-22, 8),
    to_signed(-8, 8),
    to_signed(3, 8),
    to_signed(7, 8),
    to_signed(5, 8),
    to_signed(-4, 8),
    to_signed(-16, 8),
    to_signed(-29, 8),
    to_signed(-41, 8),
    to_signed(-48, 8),
    to_signed(-48, 8),
    to_signed(-40, 8),
    to_signed(-27, 8),
    to_signed(-10, 8),
    to_signed(7, 8),
    to_signed(20, 8),
    to_signed(30, 8),
    to_signed(36, 8),
    to_signed(39, 8),
    to_signed(41, 8),
    to_signed(42, 8),
    to_signed(39, 8),
    to_signed(32, 8),
    to_signed(21, 8),
    to_signed(10, 8),
    to_signed(1, 8),
    to_signed(-3, 8),
    to_signed(-1, 8),
    to_signed(6, 8),
    to_signed(19, 8),
    to_signed(33, 8),
    to_signed(48, 8),
    to_signed(59, 8),
    to_signed(66, 8),
    to_signed(67, 8),
    to_signed(61, 8),
    to_signed(49, 8),
    to_signed(31, 8),
    to_signed(8, 8),
    to_signed(-16, 8),
    to_signed(-41, 8),
    to_signed(-64, 8),
    to_signed(-83, 8),
    to_signed(-93, 8),
    to_signed(-89, 8),
    to_signed(-71, 8),
    to_signed(-42, 8),
    to_signed(-12, 8),
    to_signed(14, 8),
    to_signed(31, 8),
    to_signed(37, 8),
    to_signed(30, 8),
    to_signed(10, 8),
    to_signed(-18, 8),
    to_signed(-46, 8),
    to_signed(-65, 8),
    to_signed(-71, 8),
    to_signed(-63, 8),
    to_signed(-45, 8),
    to_signed(-21, 8),
    to_signed(6, 8),
    to_signed(30, 8),
    to_signed(48, 8),
    to_signed(56, 8),
    to_signed(54, 8),
    to_signed(44, 8),
    to_signed(29, 8),
    to_signed(12, 8),
    to_signed(-5, 8),
    to_signed(-21, 8),
    to_signed(-33, 8),
    to_signed(-39, 8),
    to_signed(-37, 8),
    to_signed(-28, 8),
    to_signed(-15, 8),
    to_signed(-3, 8),
    to_signed(5, 8),
    to_signed(8, 8),
    to_signed(4, 8),
    to_signed(-6, 8),
    to_signed(-20, 8),
    to_signed(-34, 8),
    to_signed(-45, 8),
    to_signed(-49, 8),
    to_signed(-46, 8),
    to_signed(-38, 8),
    to_signed(-26, 8),
    to_signed(-12, 8),
    to_signed(4, 8),
    to_signed(20, 8),
    to_signed(31, 8),
    to_signed(36, 8),
    to_signed(38, 8),
    to_signed(40, 8),
    to_signed(42, 8),
    to_signed(41, 8),
    to_signed(34, 8),
    to_signed(24, 8),
    to_signed(15, 8),
    to_signed(10, 8),
    to_signed(10, 8),
    to_signed(12, 8),
    to_signed(19, 8),
    to_signed(31, 8),
    to_signed(47, 8),
    to_signed(62, 8),
    to_signed(71, 8),
    to_signed(72, 8),
    to_signed(67, 8),
    to_signed(57, 8),
    to_signed(42, 8),
    to_signed(22, 8),
    to_signed(-4, 8),
    to_signed(-31, 8),
    to_signed(-55, 8),
    to_signed(-76, 8),
    to_signed(-88, 8),
    to_signed(-90, 8),
    to_signed(-78, 8),
    to_signed(-53, 8),
    to_signed(-21, 8),
    to_signed(10, 8),
    to_signed(34, 8),
    to_signed(46, 8),
    to_signed(45, 8),
    to_signed(30, 8),
    to_signed(4, 8),
    to_signed(-27, 8),
    to_signed(-56, 8),
    to_signed(-73, 8),
    to_signed(-76, 8),
    to_signed(-64, 8),
    to_signed(-41, 8),
    to_signed(-13, 8),
    to_signed(13, 8),
    to_signed(34, 8),
    to_signed(46, 8),
    to_signed(50, 8),
    to_signed(45, 8),
    to_signed(33, 8),
    to_signed(16, 8),
    to_signed(-2, 8),
    to_signed(-18, 8),
    to_signed(-29, 8),
    to_signed(-34, 8),
    to_signed(-35, 8),
    to_signed(-30, 8),
    to_signed(-20, 8),
    to_signed(-8, 8),
    to_signed(2, 8),
    to_signed(4, 8),
    to_signed(0, 8),
    to_signed(-10, 8),
    to_signed(-21, 8),
    to_signed(-34, 8),
    to_signed(-46, 8),
    to_signed(-55, 8),
    to_signed(-58, 8),
    to_signed(-52, 8),
    to_signed(-40, 8),
    to_signed(-23, 8),
    to_signed(-5, 8),
    to_signed(12, 8),
    to_signed(26, 8),
    to_signed(36, 8),
    to_signed(43, 8),
    to_signed(48, 8),
    to_signed(50, 8),
    to_signed(50, 8),
    to_signed(45, 8),
    to_signed(37, 8),
    to_signed(27, 8),
    to_signed(20, 8),
    to_signed(17, 8),
    to_signed(16, 8),
    to_signed(17, 8),
    to_signed(23, 8),
    to_signed(33, 8),
    to_signed(46, 8),
    to_signed(57, 8),
    to_signed(63, 8),
    to_signed(65, 8),
    to_signed(63, 8),
    to_signed(56, 8),
    to_signed(42, 8),
    to_signed(21, 8),
    to_signed(-4, 8),
    to_signed(-30, 8),
    to_signed(-54, 8),
    to_signed(-75, 8),
    to_signed(-89, 8),
    to_signed(-89, 8),
    to_signed(-73, 8),
    to_signed(-44, 8),
    to_signed(-11, 8),
    to_signed(16, 8),
    to_signed(31, 8),
    to_signed(34, 8),
    to_signed(24, 8),
    to_signed(0, 8),
    to_signed(-31, 8),
    to_signed(-62, 8),
    to_signed(-81, 8),
    to_signed(-84, 8),
    to_signed(-72, 8),
    to_signed(-50, 8),
    to_signed(-21, 8),
    to_signed(10, 8),
    to_signed(36, 8),
    to_signed(53, 8),
    to_signed(58, 8),
    to_signed(54, 8),
    to_signed(43, 8),
    to_signed(28, 8),
    to_signed(10, 8),
    to_signed(-9, 8),
    to_signed(-26, 8),
    to_signed(-36, 8),
    to_signed(-39, 8),
    to_signed(-36, 8),
    to_signed(-27, 8),
    to_signed(-14, 8),
    to_signed(0, 8),
    to_signed(9, 8),
    to_signed(12, 8),
    to_signed(7, 8),
    to_signed(-3, 8),
    to_signed(-17, 8),
    to_signed(-31, 8),
    to_signed(-44, 8),
    to_signed(-51, 8),
    to_signed(-49, 8),
    to_signed(-39, 8),
    to_signed(-21, 8),
    to_signed(-1, 8),
    to_signed(18, 8),
    to_signed(34, 8),
    to_signed(44, 8),
    to_signed(50, 8),
    to_signed(52, 8),
    to_signed(53, 8),
    to_signed(51, 8),
    to_signed(45, 8),
    to_signed(36, 8),
    to_signed(26, 8),
    to_signed(20, 8),
    to_signed(17, 8),
    to_signed(18, 8),
    to_signed(20, 8),
    to_signed(25, 8),
    to_signed(35, 8),
    to_signed(48, 8),
    to_signed(60, 8),
    to_signed(67, 8),
    to_signed(67, 8),
    to_signed(64, 8),
    to_signed(58, 8),
    to_signed(46, 8),
    to_signed(27, 8),
    to_signed(1, 8),
    to_signed(-25, 8),
    to_signed(-49, 8),
    to_signed(-69, 8),
    to_signed(-87, 8),
    to_signed(-97, 8),
    to_signed(-92, 8),
    to_signed(-72, 8),
    to_signed(-41, 8),
    to_signed(-10, 8),
    to_signed(13, 8),
    to_signed(24, 8),
    to_signed(23, 8),
    to_signed(12, 8),
    to_signed(-10, 8),
    to_signed(-39, 8),
    to_signed(-63, 8),
    to_signed(-76, 8),
    to_signed(-73, 8),
    to_signed(-57, 8),
    to_signed(-34, 8),
    to_signed(-8, 8),
    to_signed(16, 8),
    to_signed(35, 8),
    to_signed(45, 8),
    to_signed(46, 8),
    to_signed(38, 8),
    to_signed(25, 8),
    to_signed(10, 8),
    to_signed(-5, 8),
    to_signed(-17, 8),
    to_signed(-25, 8),
    to_signed(-28, 8),
    to_signed(-29, 8),
    to_signed(-26, 8),
    to_signed(-18, 8),
    to_signed(-8, 8),
    to_signed(2, 8),
    to_signed(8, 8),
    to_signed(9, 8),
    to_signed(6, 8),
    to_signed(-1, 8),
    to_signed(-12, 8),
    to_signed(-26, 8),
    to_signed(-39, 8),
    to_signed(-48, 8),
    to_signed(-48, 8),
    to_signed(-39, 8),
    to_signed(-26, 8),
    to_signed(-10, 8),
    to_signed(4, 8),
    to_signed(18, 8),
    to_signed(29, 8),
    to_signed(37, 8),
    to_signed(41, 8),
    to_signed(42, 8),
    to_signed(40, 8),
    to_signed(37, 8),
    to_signed(33, 8),
    to_signed(28, 8),
    to_signed(25, 8),
    to_signed(23, 8),
    to_signed(23, 8),
    to_signed(24, 8),
    to_signed(26, 8),
    to_signed(30, 8),
    to_signed(37, 8),
    to_signed(43, 8),
    to_signed(46, 8),
    to_signed(47, 8),
    to_signed(47, 8),
    to_signed(45, 8),
    to_signed(38, 8),
    to_signed(25, 8),
    to_signed(6, 8),
    to_signed(-15, 8),
    to_signed(-38, 8),
    to_signed(-60, 8),
    to_signed(-80, 8),
    to_signed(-91, 8),
    to_signed(-87, 8),
    to_signed(-67, 8),
    to_signed(-39, 8),
    to_signed(-10, 8),
    to_signed(13, 8),
    to_signed(26, 8),
    to_signed(29, 8),
    to_signed(20, 8),
    to_signed(-2, 8),
    to_signed(-29, 8),
    to_signed(-54, 8),
    to_signed(-68, 8),
    to_signed(-68, 8),
    to_signed(-56, 8),
    to_signed(-35, 8),
    to_signed(-10, 8),
    to_signed(16, 8),
    to_signed(38, 8),
    to_signed(50, 8),
    to_signed(52, 8),
    to_signed(46, 8),
    to_signed(34, 8),
    to_signed(20, 8),
    to_signed(7, 8),
    to_signed(-3, 8),
    to_signed(-11, 8),
    to_signed(-17, 8),
    to_signed(-20, 8),
    to_signed(-18, 8),
    to_signed(-12, 8),
    to_signed(-4, 8),
    to_signed(2, 8),
    to_signed(6, 8),
    to_signed(5, 8),
    to_signed(1, 8),
    to_signed(-5, 8),
    to_signed(-16, 8),
    to_signed(-32, 8),
    to_signed(-49, 8),
    to_signed(-58, 8),
    to_signed(-55, 8),
    to_signed(-43, 8),
    to_signed(-26, 8),
    to_signed(-8, 8),
    to_signed(9, 8),
    to_signed(25, 8),
    to_signed(38, 8),
    to_signed(46, 8),
    to_signed(49, 8),
    to_signed(48, 8),
    to_signed(45, 8),
    to_signed(40, 8),
    to_signed(34, 8),
    to_signed(26, 8),
    to_signed(21, 8),
    to_signed(19, 8),
    to_signed(21, 8),
    to_signed(25, 8),
    to_signed(29, 8),
    to_signed(35, 8),
    to_signed(42, 8),
    to_signed(49, 8),
    to_signed(55, 8),
    to_signed(59, 8),
    to_signed(60, 8),
    to_signed(56, 8),
    to_signed(47, 8),
    to_signed(32, 8),
    to_signed(12, 8),
    to_signed(-12, 8),
    to_signed(-37, 8),
    to_signed(-61, 8),
    to_signed(-80, 8),
    to_signed(-88, 8),
    to_signed(-80, 8),
    to_signed(-57, 8),
    to_signed(-27, 8),
    to_signed(1, 8),
    to_signed(22, 8),
    to_signed(32, 8),
    to_signed(29, 8),
    to_signed(14, 8),
    to_signed(-11, 8),
    to_signed(-38, 8),
    to_signed(-61, 8),
    to_signed(-72, 8),
    to_signed(-69, 8),
    to_signed(-53, 8),
    to_signed(-29, 8),
    to_signed(-1, 8),
    to_signed(25, 8),
    to_signed(45, 8),
    to_signed(54, 8),
    to_signed(53, 8),
    to_signed(46, 8),
    to_signed(34, 8),
    to_signed(18, 8),
    to_signed(2, 8),
    to_signed(-13, 8),
    to_signed(-25, 8),
    to_signed(-33, 8),
    to_signed(-35, 8),
    to_signed(-30, 8),
    to_signed(-21, 8),
    to_signed(-9, 8),
    to_signed(2, 8),
    to_signed(10, 8),
    to_signed(13, 8),
    to_signed(9, 8),
    to_signed(-1, 8),
    to_signed(-19, 8),
    to_signed(-41, 8),
    to_signed(-60, 8),
    to_signed(-67, 8),
    to_signed(-62, 8),
    to_signed(-46, 8),
    to_signed(-25, 8),
    to_signed(-3, 8),
    to_signed(18, 8),
    to_signed(36, 8),
    to_signed(49, 8),
    to_signed(54, 8),
    to_signed(54, 8),
    to_signed(50, 8),
    to_signed(44, 8),
    to_signed(36, 8),
    to_signed(26, 8),
    to_signed(17, 8),
    to_signed(11, 8),
    to_signed(11, 8),
    to_signed(15, 8),
    to_signed(20, 8),
    to_signed(28, 8),
    to_signed(38, 8),
    to_signed(49, 8),
    to_signed(58, 8),
    to_signed(63, 8),
    to_signed(63, 8),
    to_signed(58, 8),
    to_signed(49, 8),
    to_signed(35, 8),
    to_signed(15, 8),
    to_signed(-10, 8),
    to_signed(-37, 8),
    to_signed(-63, 8),
    to_signed(-84, 8),
    to_signed(-96, 8),
    to_signed(-95, 8),
    to_signed(-79, 8),
    to_signed(-51, 8),
    to_signed(-19, 8),
    to_signed(10, 8),
    to_signed(29, 8),
    to_signed(35, 8),
    to_signed(27, 8),
    to_signed(8, 8),
    to_signed(-18, 8),
    to_signed(-45, 8),
    to_signed(-65, 8),
    to_signed(-71, 8),
    to_signed(-63, 8),
    to_signed(-44, 8),
    to_signed(-19, 8),
    to_signed(8, 8),
    to_signed(29, 8),
    to_signed(41, 8),
    to_signed(42, 8),
    to_signed(35, 8),
    to_signed(23, 8),
    to_signed(6, 8),
    to_signed(-13, 8),
    to_signed(-29, 8),
    to_signed(-39, 8),
    to_signed(-43, 8),
    to_signed(-41, 8),
    to_signed(-35, 8),
    to_signed(-24, 8),
    to_signed(-11, 8),
    to_signed(3, 8),
    to_signed(17, 8),
    to_signed(24, 8),
    to_signed(22, 8),
    to_signed(11, 8),
    to_signed(-5, 8),
    to_signed(-25, 8),
    to_signed(-46, 8),
    to_signed(-63, 8),
    to_signed(-69, 8),
    to_signed(-62, 8),
    to_signed(-43, 8),
    to_signed(-17, 8),
    to_signed(10, 8),
    to_signed(34, 8),
    to_signed(52, 8),
    to_signed(63, 8),
    to_signed(67, 8),
    to_signed(63, 8),
    to_signed(51, 8),
    to_signed(36, 8),
    to_signed(23, 8),
    to_signed(13, 8),
    to_signed(8, 8),
    to_signed(9, 8),
    to_signed(14, 8),
    to_signed(21, 8),
    to_signed(30, 8),
    to_signed(40, 8),
    to_signed(48, 8),
    to_signed(52, 8),
    to_signed(52, 8),
    to_signed(48, 8),
    to_signed(45, 8),
    to_signed(40, 8),
    to_signed(33, 8),
    to_signed(22, 8),
    to_signed(6, 8),
    to_signed(-12, 8),
    to_signed(-31, 8),
    to_signed(-51, 8),
    to_signed(-71, 8),
    to_signed(-86, 8),
    to_signed(-89, 8),
    to_signed(-77, 8),
    to_signed(-51, 8),
    to_signed(-22, 8),
    to_signed(3, 8),
    to_signed(19, 8),
    to_signed(25, 8),
    to_signed(18, 8),
    to_signed(0, 8),
    to_signed(-26, 8),
    to_signed(-53, 8),
    to_signed(-72, 8),
    to_signed(-77, 8),
    to_signed(-67, 8),
    to_signed(-48, 8),
    to_signed(-22, 8),
    to_signed(6, 8),
    to_signed(31, 8),
    to_signed(48, 8),
    to_signed(51, 8),
    to_signed(43, 8),
    to_signed(29, 8),
    to_signed(14, 8),
    to_signed(2, 8),
    to_signed(-8, 8),
    to_signed(-16, 8),
    to_signed(-20, 8),
    to_signed(-19, 8),
    to_signed(-12, 8),
    to_signed(-2, 8),
    to_signed(8, 8),
    to_signed(18, 8),
    to_signed(25, 8),
    to_signed(27, 8),
    to_signed(24, 8),
    to_signed(15, 8),
    to_signed(0, 8),
    to_signed(-19, 8),
    to_signed(-37, 8),
    to_signed(-51, 8),
    to_signed(-54, 8),
    to_signed(-47, 8),
    to_signed(-30, 8),
    to_signed(-6, 8),
    to_signed(19, 8),
    to_signed(41, 8),
    to_signed(57, 8),
    to_signed(66, 8),
    to_signed(66, 8),
    to_signed(59, 8),
    to_signed(47, 8),
    to_signed(34, 8),
    to_signed(22, 8),
    to_signed(10, 8),
    to_signed(2, 8),
    to_signed(-1, 8),
    to_signed(3, 8),
    to_signed(9, 8),
    to_signed(17, 8),
    to_signed(25, 8),
    to_signed(33, 8),
    to_signed(39, 8),
    to_signed(43, 8),
    to_signed(43, 8),
    to_signed(40, 8),
    to_signed(37, 8),
    to_signed(34, 8),
    to_signed(28, 8),
    to_signed(17, 8),
    to_signed(2, 8),
    to_signed(-15, 8),
    to_signed(-33, 8),
    to_signed(-52, 8),
    to_signed(-72, 8),
    to_signed(-85, 8),
    to_signed(-84, 8),
    to_signed(-68, 8),
    to_signed(-42, 8),
    to_signed(-14, 8),
    to_signed(9, 8),
    to_signed(23, 8),
    to_signed(27, 8),
    to_signed(21, 8),
    to_signed(4, 8),
    to_signed(-21, 8),
    to_signed(-45, 8),
    to_signed(-58, 8),
    to_signed(-57, 8),
    to_signed(-44, 8),
    to_signed(-22, 8),
    to_signed(4, 8),
    to_signed(29, 8),
    to_signed(46, 8),
    to_signed(55, 8),
    to_signed(54, 8),
    to_signed(47, 8),
    to_signed(36, 8),
    to_signed(23, 8),
    to_signed(9, 8),
    to_signed(-3, 8),
    to_signed(-9, 8),
    to_signed(-12, 8),
    to_signed(-12, 8),
    to_signed(-10, 8),
    to_signed(-4, 8),
    to_signed(5, 8),
    to_signed(15, 8),
    to_signed(22, 8),
    to_signed(23, 8),
    to_signed(20, 8),
    to_signed(11, 8),
    to_signed(-4, 8),
    to_signed(-23, 8),
    to_signed(-41, 8),
    to_signed(-53, 8),
    to_signed(-53, 8),
    to_signed(-43, 8),
    to_signed(-28, 8),
    to_signed(-11, 8),
    to_signed(7, 8),
    to_signed(23, 8),
    to_signed(37, 8),
    to_signed(42, 8),
    to_signed(38, 8),
    to_signed(30, 8),
    to_signed(23, 8),
    to_signed(17, 8),
    to_signed(10, 8),
    to_signed(3, 8),
    to_signed(-3, 8),
    to_signed(-5, 8),
    to_signed(-2, 8),
    to_signed(2, 8),
    to_signed(6, 8),
    to_signed(13, 8),
    to_signed(22, 8),
    to_signed(31, 8),
    to_signed(38, 8),
    to_signed(42, 8),
    to_signed(43, 8),
    to_signed(40, 8),
    to_signed(34, 8),
    to_signed(21, 8),
    to_signed(3, 8),
    to_signed(-18, 8),
    to_signed(-41, 8),
    to_signed(-65, 8),
    to_signed(-84, 8),
    to_signed(-94, 8),
    to_signed(-88, 8),
    to_signed(-66, 8),
    to_signed(-36, 8),
    to_signed(-5, 8),
    to_signed(20, 8),
    to_signed(37, 8),
    to_signed(44, 8),
    to_signed(37, 8),
    to_signed(16, 8),
    to_signed(-12, 8),
    to_signed(-36, 8),
    to_signed(-50, 8),
    to_signed(-50, 8),
    to_signed(-40, 8),
    to_signed(-21, 8),
    to_signed(2, 8),
    to_signed(26, 8),
    to_signed(43, 8),
    to_signed(51, 8),
    to_signed(49, 8),
    to_signed(41, 8),
    to_signed(30, 8),
    to_signed(17, 8),
    to_signed(4, 8),
    to_signed(-8, 8),
    to_signed(-17, 8),
    to_signed(-21, 8),
    to_signed(-23, 8),
    to_signed(-23, 8),
    to_signed(-19, 8),
    to_signed(-11, 8),
    to_signed(0, 8),
    to_signed(9, 8),
    to_signed(13, 8),
    to_signed(10, 8),
    to_signed(1, 8),
    to_signed(-17, 8),
    to_signed(-40, 8),
    to_signed(-63, 8),
    to_signed(-79, 8),
    to_signed(-83, 8),
    to_signed(-75, 8),
    to_signed(-58, 8),
    to_signed(-34, 8),
    to_signed(-9, 8),
    to_signed(16, 8),
    to_signed(34, 8),
    to_signed(41, 8),
    to_signed(39, 8),
    to_signed(32, 8),
    to_signed(24, 8),
    to_signed(16, 8),
    to_signed(6, 8),
    to_signed(-3, 8),
    to_signed(-7, 8),
    to_signed(-5, 8),
    to_signed(0, 8),
    to_signed(5, 8),
    to_signed(11, 8),
    to_signed(20, 8),
    to_signed(32, 8),
    to_signed(43, 8),
    to_signed(50, 8),
    to_signed(51, 8),
    to_signed(50, 8),
    to_signed(47, 8),
    to_signed(39, 8),
    to_signed(24, 8),
    to_signed(4, 8),
    to_signed(-17, 8),
    to_signed(-34, 8),
    to_signed(-49, 8),
    to_signed(-61, 8),
    to_signed(-67, 8),
    to_signed(-62, 8),
    to_signed(-44, 8),
    to_signed(-19, 8),
    to_signed(5, 8),
    to_signed(25, 8),
    to_signed(36, 8),
    to_signed(37, 8),
    to_signed(25, 8),
    to_signed(3, 8),
    to_signed(-24, 8),
    to_signed(-47, 8),
    to_signed(-59, 8),
    to_signed(-57, 8),
    to_signed(-44, 8),
    to_signed(-22, 8),
    to_signed(3, 8),
    to_signed(27, 8),
    to_signed(43, 8),
    to_signed(48, 8),
    to_signed(44, 8),
    to_signed(35, 8),
    to_signed(23, 8),
    to_signed(9, 8),
    to_signed(-4, 8),
    to_signed(-15, 8),
    to_signed(-21, 8),
    to_signed(-23, 8),
    to_signed(-23, 8),
    to_signed(-23, 8),
    to_signed(-21, 8),
    to_signed(-16, 8),
    to_signed(-9, 8),
    to_signed(-3, 8),
    to_signed(-1, 8),
    to_signed(-4, 8),
    to_signed(-12, 8),
    to_signed(-25, 8),
    to_signed(-43, 8),
    to_signed(-61, 8),
    to_signed(-73, 8),
    to_signed(-73, 8),
    to_signed(-62, 8),
    to_signed(-42, 8),
    to_signed(-19, 8),
    to_signed(6, 8),
    to_signed(29, 8),
    to_signed(44, 8),
    to_signed(50, 8),
    to_signed(47, 8),
    to_signed(40, 8),
    to_signed(32, 8),
    to_signed(24, 8),
    to_signed(16, 8),
    to_signed(10, 8),
    to_signed(7, 8),
    to_signed(9, 8),
    to_signed(12, 8),
    to_signed(17, 8),
    to_signed(24, 8),
    to_signed(34, 8),
    to_signed(47, 8),
    to_signed(58, 8),
    to_signed(66, 8),
    to_signed(69, 8),
    to_signed(69, 8),
    to_signed(66, 8),
    to_signed(59, 8),
    to_signed(46, 8),
    to_signed(29, 8),
    to_signed(11, 8),
    to_signed(-6, 8),
    to_signed(-26, 8),
    to_signed(-46, 8),
    to_signed(-63, 8),
    to_signed(-67, 8),
    to_signed(-58, 8),
    to_signed(-39, 8),
    to_signed(-16, 8),
    to_signed(5, 8),
    to_signed(21, 8),
    to_signed(30, 8),
    to_signed(28, 8),
    to_signed(15, 8),
    to_signed(-8, 8),
    to_signed(-33, 8),
    to_signed(-51, 8),
    to_signed(-57, 8),
    to_signed(-50, 8),
    to_signed(-32, 8),
    to_signed(-8, 8),
    to_signed(14, 8),
    to_signed(29, 8),
    to_signed(36, 8),
    to_signed(36, 8),
    to_signed(31, 8),
    to_signed(22, 8),
    to_signed(10, 8),
    to_signed(-3, 8),
    to_signed(-13, 8),
    to_signed(-21, 8),
    to_signed(-24, 8),
    to_signed(-26, 8),
    to_signed(-28, 8),
    to_signed(-28, 8),
    to_signed(-22, 8),
    to_signed(-13, 8),
    to_signed(-4, 8),
    to_signed(1, 8),
    to_signed(3, 8),
    to_signed(1, 8),
    to_signed(-6, 8),
    to_signed(-20, 8),
    to_signed(-37, 8),
    to_signed(-53, 8),
    to_signed(-59, 8),
    to_signed(-54, 8),
    to_signed(-40, 8),
    to_signed(-22, 8),
    to_signed(-3, 8),
    to_signed(15, 8),
    to_signed(31, 8),
    to_signed(42, 8),
    to_signed(46, 8),
    to_signed(44, 8),
    to_signed(40, 8),
    to_signed(34, 8),
    to_signed(27, 8),
    to_signed(21, 8),
    to_signed(18, 8),
    to_signed(19, 8),
    to_signed(22, 8),
    to_signed(26, 8),
    to_signed(32, 8),
    to_signed(37, 8),
    to_signed(43, 8),
    to_signed(48, 8),
    to_signed(54, 8),
    to_signed(58, 8),
    to_signed(60, 8),
    to_signed(59, 8),
    to_signed(50, 8),
    to_signed(34, 8),
    to_signed(13, 8),
    to_signed(-8, 8),
    to_signed(-29, 8),
    to_signed(-52, 8),
    to_signed(-76, 8),
    to_signed(-91, 8),
    to_signed(-92, 8),
    to_signed(-76, 8),
    to_signed(-50, 8),
    to_signed(-21, 8),
    to_signed(3, 8),
    to_signed(21, 8),
    to_signed(29, 8),
    to_signed(24, 8),
    to_signed(5, 8),
    to_signed(-24, 8),
    to_signed(-51, 8),
    to_signed(-66, 8),
    to_signed(-68, 8),
    to_signed(-59, 8),
    to_signed(-42, 8),
    to_signed(-21, 8),
    to_signed(1, 8),
    to_signed(18, 8),
    to_signed(29, 8),
    to_signed(33, 8),
    to_signed(31, 8),
    to_signed(27, 8),
    to_signed(21, 8),
    to_signed(12, 8),
    to_signed(2, 8),
    to_signed(-9, 8),
    to_signed(-18, 8),
    to_signed(-24, 8),
    to_signed(-26, 8),
    to_signed(-24, 8),
    to_signed(-15, 8),
    to_signed(-4, 8),
    to_signed(6, 8),
    to_signed(11, 8),
    to_signed(10, 8),
    to_signed(4, 8),
    to_signed(-8, 8),
    to_signed(-25, 8),
    to_signed(-44, 8),
    to_signed(-58, 8),
    to_signed(-64, 8),
    to_signed(-58, 8),
    to_signed(-43, 8),
    to_signed(-23, 8),
    to_signed(-2, 8),
    to_signed(18, 8),
    to_signed(35, 8),
    to_signed(47, 8),
    to_signed(52, 8),
    to_signed(52, 8),
    to_signed(49, 8),
    to_signed(42, 8),
    to_signed(31, 8),
    to_signed(20, 8),
    to_signed(12, 8),
    to_signed(8, 8),
    to_signed(7, 8),
    to_signed(8, 8),
    to_signed(12, 8),
    to_signed(21, 8),
    to_signed(33, 8),
    to_signed(46, 8),
    to_signed(54, 8),
    to_signed(58, 8),
    to_signed(58, 8),
    to_signed(53, 8),
    to_signed(41, 8),
    to_signed(21, 8),
    to_signed(-1, 8),
    to_signed(-22, 8),
    to_signed(-39, 8),
    to_signed(-58, 8),
    to_signed(-76, 8),
    to_signed(-89, 8),
    to_signed(-89, 8),
    to_signed(-73, 8),
    to_signed(-47, 8),
    to_signed(-21, 8),
    to_signed(-1, 8),
    to_signed(12, 8),
    to_signed(17, 8),
    to_signed(11, 8),
    to_signed(-7, 8),
    to_signed(-33, 8),
    to_signed(-55, 8),
    to_signed(-65, 8),
    to_signed(-62, 8),
    to_signed(-48, 8),
    to_signed(-29, 8),
    to_signed(-6, 8),
    to_signed(16, 8),
    to_signed(34, 8),
    to_signed(44, 8),
    to_signed(44, 8),
    to_signed(39, 8),
    to_signed(31, 8),
    to_signed(23, 8),
    to_signed(14, 8),
    to_signed(5, 8),
    to_signed(-5, 8),
    to_signed(-13, 8),
    to_signed(-20, 8),
    to_signed(-22, 8),
    to_signed(-19, 8),
    to_signed(-11, 8),
    to_signed(0, 8),
    to_signed(9, 8),
    to_signed(14, 8),
    to_signed(15, 8),
    to_signed(10, 8),
    to_signed(-2, 8),
    to_signed(-19, 8),
    to_signed(-36, 8),
    to_signed(-47, 8),
    to_signed(-47, 8),
    to_signed(-39, 8),
    to_signed(-24, 8),
    to_signed(-6, 8),
    to_signed(12, 8),
    to_signed(30, 8),
    to_signed(44, 8),
    to_signed(50, 8),
    to_signed(50, 8),
    to_signed(47, 8),
    to_signed(43, 8),
    to_signed(37, 8),
    to_signed(28, 8),
    to_signed(20, 8),
    to_signed(14, 8),
    to_signed(12, 8),
    to_signed(12, 8),
    to_signed(13, 8),
    to_signed(16, 8),
    to_signed(22, 8),
    to_signed(32, 8),
    to_signed(43, 8),
    to_signed(51, 8),
    to_signed(54, 8),
    to_signed(52, 8),
    to_signed(47, 8),
    to_signed(35, 8),
    to_signed(17, 8),
    to_signed(-3, 8),
    to_signed(-22, 8),
    to_signed(-39, 8),
    to_signed(-56, 8),
    to_signed(-74, 8),
    to_signed(-86, 8),
    to_signed(-86, 8),
    to_signed(-71, 8),
    to_signed(-46, 8),
    to_signed(-20, 8),
    to_signed(1, 8),
    to_signed(16, 8),
    to_signed(21, 8),
    to_signed(16, 8),
    to_signed(0, 8),
    to_signed(-23, 8),
    to_signed(-43, 8),
    to_signed(-53, 8),
    to_signed(-51, 8),
    to_signed(-40, 8),
    to_signed(-22, 8),
    to_signed(0, 8),
    to_signed(20, 8),
    to_signed(36, 8),
    to_signed(44, 8),
    to_signed(44, 8),
    to_signed(39, 8),
    to_signed(31, 8),
    to_signed(23, 8),
    to_signed(15, 8),
    to_signed(6, 8),
    to_signed(-2, 8),
    to_signed(-9, 8),
    to_signed(-15, 8),
    to_signed(-18, 8),
    to_signed(-15, 8),
    to_signed(-6, 8),
    to_signed(4, 8),
    to_signed(11, 8),
    to_signed(15, 8),
    to_signed(15, 8),
    to_signed(11, 8),
    to_signed(0, 8),
    to_signed(-17, 8),
    to_signed(-35, 8),
    to_signed(-48, 8),
    to_signed(-52, 8),
    to_signed(-47, 8),
    to_signed(-35, 8),
    to_signed(-20, 8),
    to_signed(-3, 8),
    to_signed(13, 8),
    to_signed(26, 8),
    to_signed(31, 8),
    to_signed(30, 8),
    to_signed(26, 8),
    to_signed(22, 8),
    to_signed(16, 8),
    to_signed(10, 8),
    to_signed(5, 8),
    to_signed(3, 8),
    to_signed(4, 8),
    to_signed(8, 8),
    to_signed(12, 8),
    to_signed(17, 8),
    to_signed(24, 8),
    to_signed(34, 8),
    to_signed(42, 8),
    to_signed(47, 8),
    to_signed(48, 8),
    to_signed(47, 8),
    to_signed(44, 8),
    to_signed(35, 8),
    to_signed(20, 8),
    to_signed(0, 8),
    to_signed(-22, 8),
    to_signed(-44, 8),
    to_signed(-66, 8),
    to_signed(-82, 8),
    to_signed(-88, 8),
    to_signed(-77, 8),
    to_signed(-53, 8),
    to_signed(-23, 8),
    to_signed(4, 8),
    to_signed(23, 8),
    to_signed(33, 8),
    to_signed(31, 8),
    to_signed(17, 8),
    to_signed(-6, 8),
    to_signed(-32, 8),
    to_signed(-51, 8),
    to_signed(-58, 8),
    to_signed(-52, 8),
    to_signed(-37, 8),
    to_signed(-16, 8),
    to_signed(7, 8),
    to_signed(26, 8),
    to_signed(39, 8),
    to_signed(43, 8),
    to_signed(41, 8),
    to_signed(35, 8),
    to_signed(27, 8),
    to_signed(17, 8),
    to_signed(5, 8),
    to_signed(-7, 8),
    to_signed(-15, 8),
    to_signed(-20, 8),
    to_signed(-21, 8),
    to_signed(-20, 8),
    to_signed(-16, 8),
    to_signed(-9, 8),
    to_signed(-3, 8),
    to_signed(0, 8),
    to_signed(1, 8),
    to_signed(-3, 8),
    to_signed(-10, 8),
    to_signed(-23, 8),
    to_signed(-41, 8),
    to_signed(-57, 8),
    to_signed(-66, 8),
    to_signed(-63, 8),
    to_signed(-50, 8),
    to_signed(-31, 8),
    to_signed(-12, 8),
    to_signed(7, 8),
    to_signed(23, 8),
    to_signed(36, 8),
    to_signed(43, 8),
    to_signed(46, 8),
    to_signed(45, 8),
    to_signed(39, 8),
    to_signed(30, 8),
    to_signed(20, 8),
    to_signed(11, 8),
    to_signed(6, 8),
    to_signed(6, 8),
    to_signed(9, 8),
    to_signed(15, 8),
    to_signed(25, 8),
    to_signed(39, 8),
    to_signed(52, 8),
    to_signed(61, 8),
    to_signed(64, 8),
    to_signed(61, 8),
    to_signed(56, 8),
    to_signed(47, 8),
    to_signed(32, 8),
    to_signed(11, 8),
    to_signed(-12, 8),
    to_signed(-34, 8),
    to_signed(-53, 8),
    to_signed(-71, 8),
    to_signed(-83, 8),
    to_signed(-82, 8),
    to_signed(-64, 8),
    to_signed(-35, 8),
    to_signed(-4, 8),
    to_signed(19, 8),
    to_signed(32, 8),
    to_signed(34, 8),
    to_signed(25, 8),
    to_signed(5, 8),
    to_signed(-24, 8),
    to_signed(-52, 8),
    to_signed(-69, 8),
    to_signed(-69, 8),
    to_signed(-55, 8),
    to_signed(-33, 8),
    to_signed(-7, 8),
    to_signed(18, 8),
    to_signed(38, 8),
    to_signed(50, 8),
    to_signed(52, 8),
    to_signed(45, 8),
    to_signed(33, 8),
    to_signed(18, 8),
    to_signed(1, 8),
    to_signed(-15, 8),
    to_signed(-28, 8),
    to_signed(-35, 8),
    to_signed(-35, 8),
    to_signed(-30, 8),
    to_signed(-22, 8),
    to_signed(-11, 8),
    to_signed(0, 8),
    to_signed(9, 8),
    to_signed(13, 8),
    to_signed(11, 8),
    to_signed(5, 8),
    to_signed(-5, 8),
    to_signed(-19, 8),
    to_signed(-35, 8),
    to_signed(-46, 8),
    to_signed(-48, 8),
    to_signed(-39, 8),
    to_signed(-22, 8),
    to_signed(-3, 8),
    to_signed(16, 8),
    to_signed(34, 8),
    to_signed(48, 8),
    to_signed(56, 8),
    to_signed(56, 8),
    to_signed(50, 8),
    to_signed(42, 8),
    to_signed(34, 8),
    to_signed(26, 8),
    to_signed(17, 8),
    to_signed(12, 8),
    to_signed(10, 8),
    to_signed(13, 8),
    to_signed(17, 8),
    to_signed(25, 8),
    to_signed(37, 8),
    to_signed(50, 8),
    to_signed(61, 8),
    to_signed(65, 8),
    to_signed(60, 8),
    to_signed(51, 8),
    to_signed(41, 8),
    to_signed(30, 8),
    to_signed(15, 8),
    to_signed(-2, 8),
    to_signed(-20, 8),
    to_signed(-37, 8),
    to_signed(-55, 8),
    to_signed(-73, 8),
    to_signed(-86, 8),
    to_signed(-85, 8),
    to_signed(-69, 8),
    to_signed(-42, 8),
    to_signed(-14, 8),
    to_signed(9, 8),
    to_signed(23, 8),
    to_signed(27, 8),
    to_signed(20, 8),
    to_signed(1, 8),
    to_signed(-27, 8),
    to_signed(-52, 8),
    to_signed(-66, 8),
    to_signed(-65, 8),
    to_signed(-53, 8),
    to_signed(-33, 8),
    to_signed(-10, 8),
    to_signed(14, 8),
    to_signed(33, 8),
    to_signed(43, 8),
    to_signed(43, 8),
    to_signed(35, 8),
    to_signed(24, 8),
    to_signed(11, 8),
    to_signed(-2, 8),
    to_signed(-13, 8),
    to_signed(-20, 8),
    to_signed(-23, 8),
    to_signed(-21, 8),
    to_signed(-17, 8),
    to_signed(-10, 8),
    to_signed(-2, 8),
    to_signed(7, 8),
    to_signed(13, 8),
    to_signed(16, 8),
    to_signed(15, 8),
    to_signed(11, 8),
    to_signed(2, 8),
    to_signed(-13, 8),
    to_signed(-29, 8),
    to_signed(-40, 8),
    to_signed(-42, 8),
    to_signed(-34, 8),
    to_signed(-19, 8),
    to_signed(0, 8),
    to_signed(19, 8),
    to_signed(35, 8),
    to_signed(47, 8),
    to_signed(52, 8),
    to_signed(50, 8),
    to_signed(43, 8),
    to_signed(36, 8),
    to_signed(27, 8),
    to_signed(17, 8),
    to_signed(9, 8),
    to_signed(5, 8),
    to_signed(6, 8),
    to_signed(11, 8),
    to_signed(16, 8),
    to_signed(23, 8),
    to_signed(30, 8),
    to_signed(38, 8),
    to_signed(44, 8),
    to_signed(46, 8),
    to_signed(44, 8),
    to_signed(40, 8),
    to_signed(35, 8),
    to_signed(27, 8),
    to_signed(12, 8),
    to_signed(-8, 8),
    to_signed(-30, 8),
    to_signed(-51, 8),
    to_signed(-71, 8),
    to_signed(-87, 8),
    to_signed(-94, 8),
    to_signed(-85, 8),
    to_signed(-63, 8),
    to_signed(-33, 8),
    to_signed(-6, 8),
    to_signed(14, 8),
    to_signed(24, 8),
    to_signed(23, 8),
    to_signed(12, 8),
    to_signed(-9, 8),
    to_signed(-34, 8),
    to_signed(-53, 8),
    to_signed(-60, 8),
    to_signed(-55, 8),
    to_signed(-40, 8),
    to_signed(-19, 8),
    to_signed(3, 8),
    to_signed(24, 8),
    to_signed(38, 8),
    to_signed(44, 8),
    to_signed(41, 8),
    to_signed(34, 8),
    to_signed(23, 8),
    to_signed(12, 8),
    to_signed(0, 8),
    to_signed(-11, 8),
    to_signed(-19, 8),
    to_signed(-22, 8),
    to_signed(-20, 8),
    to_signed(-14, 8),
    to_signed(-6, 8),
    to_signed(4, 8),
    to_signed(12, 8),
    to_signed(17, 8),
    to_signed(17, 8),
    to_signed(11, 8),
    to_signed(0, 8),
    to_signed(-16, 8),
    to_signed(-33, 8),
    to_signed(-46, 8),
    to_signed(-51, 8),
    to_signed(-48, 8),
    to_signed(-37, 8),
    to_signed(-20, 8),
    to_signed(-2, 8),
    to_signed(16, 8),
    to_signed(32, 8),
    to_signed(43, 8),
    to_signed(48, 8),
    to_signed(47, 8),
    to_signed(41, 8),
    to_signed(31, 8),
    to_signed(18, 8),
    to_signed(6, 8),
    to_signed(-4, 8),
    to_signed(-8, 8),
    to_signed(-7, 8),
    to_signed(-3, 8),
    to_signed(5, 8),
    to_signed(16, 8),
    to_signed(30, 8),
    to_signed(43, 8),
    to_signed(51, 8),
    to_signed(53, 8),
    to_signed(48, 8),
    to_signed(40, 8),
    to_signed(30, 8),
    to_signed(16, 8),
    to_signed(-2, 8),
    to_signed(-23, 8),
    to_signed(-45, 8),
    to_signed(-66, 8),
    to_signed(-82, 8),
    to_signed(-90, 8),
    to_signed(-85, 8),
    to_signed(-67, 8),
    to_signed(-40, 8),
    to_signed(-11, 8),
    to_signed(13, 8),
    to_signed(26, 8),
    to_signed(27, 8),
    to_signed(16, 8),
    to_signed(-4, 8),
    to_signed(-30, 8),
    to_signed(-53, 8),
    to_signed(-66, 8),
    to_signed(-64, 8),
    to_signed(-50, 8),
    to_signed(-28, 8),
    to_signed(-3, 8),
    to_signed(21, 8),
    to_signed(38, 8),
    to_signed(46, 8),
    to_signed(46, 8),
    to_signed(39, 8),
    to_signed(28, 8),
    to_signed(15, 8),
    to_signed(1, 8),
    to_signed(-14, 8),
    to_signed(-26, 8),
    to_signed(-33, 8),
    to_signed(-32, 8),
    to_signed(-26, 8),
    to_signed(-16, 8),
    to_signed(-5, 8),
    to_signed(6, 8),
    to_signed(14, 8),
    to_signed(18, 8),
    to_signed(15, 8),
    to_signed(6, 8),
    to_signed(-8, 8),
    to_signed(-25, 8),
    to_signed(-41, 8),
    to_signed(-52, 8),
    to_signed(-54, 8),
    to_signed(-46, 8),
    to_signed(-30, 8),
    to_signed(-9, 8),
    to_signed(12, 8),
    to_signed(30, 8),
    to_signed(42, 8),
    to_signed(49, 8),
    to_signed(52, 8),
    to_signed(51, 8),
    to_signed(46, 8),
    to_signed(38, 8),
    to_signed(26, 8),
    to_signed(14, 8),
    to_signed(5, 8),
    to_signed(1, 8),
    to_signed(0, 8),
    to_signed(5, 8),
    to_signed(15, 8),
    to_signed(31, 8),
    to_signed(48, 8),
    to_signed(61, 8),
    to_signed(68, 8),
    to_signed(67, 8),
    to_signed(61, 8),
    to_signed(52, 8),
    to_signed(39, 8),
    to_signed(20, 8),
    to_signed(-1, 8),
    to_signed(-23, 8),
    to_signed(-43, 8),
    to_signed(-61, 8),
    to_signed(-76, 8),
    to_signed(-83, 8),
    to_signed(-77, 8),
    to_signed(-57, 8),
    to_signed(-30, 8),
    to_signed(-2, 8),
    to_signed(21, 8),
    to_signed(34, 8),
    to_signed(34, 8),
    to_signed(23, 8),
    to_signed(2, 8),
    to_signed(-25, 8),
    to_signed(-47, 8),
    to_signed(-58, 8),
    to_signed(-55, 8),
    to_signed(-41, 8),
    to_signed(-20, 8),
    to_signed(5, 8),
    to_signed(27, 8),
    to_signed(43, 8),
    to_signed(49, 8),
    to_signed(48, 8),
    to_signed(40, 8),
    to_signed(28, 8),
    to_signed(14, 8),
    to_signed(0, 8),
    to_signed(-14, 8),
    to_signed(-24, 8),
    to_signed(-30, 8),
    to_signed(-29, 8),
    to_signed(-23, 8),
    to_signed(-13, 8),
    to_signed(0, 8),
    to_signed(12, 8),
    to_signed(20, 8),
    to_signed(23, 8),
    to_signed(20, 8),
    to_signed(11, 8),
    to_signed(-3, 8),
    to_signed(-21, 8),
    to_signed(-36, 8),
    to_signed(-45, 8),
    to_signed(-45, 8),
    to_signed(-36, 8),
    to_signed(-21, 8),
    to_signed(-2, 8),
    to_signed(17, 8),
    to_signed(34, 8),
    to_signed(47, 8),
    to_signed(53, 8),
    to_signed(55, 8),
    to_signed(53, 8),
    to_signed(48, 8),
    to_signed(39, 8),
    to_signed(26, 8),
    to_signed(12, 8),
    to_signed(2, 8),
    to_signed(-3, 8),
    to_signed(-4, 8),
    to_signed(-1, 8),
    to_signed(8, 8),
    to_signed(21, 8),
    to_signed(36, 8),
    to_signed(47, 8),
    to_signed(54, 8),
    to_signed(54, 8),
    to_signed(50, 8),
    to_signed(42, 8),
    to_signed(29, 8),
    to_signed(10, 8),
    to_signed(-10, 8),
    to_signed(-30, 8),
    to_signed(-51, 8),
    to_signed(-74, 8),
    to_signed(-94, 8),
    to_signed(-104, 8),
    to_signed(-98, 8),
    to_signed(-76, 8),
    to_signed(-47, 8),
    to_signed(-17, 8),
    to_signed(8, 8),
    to_signed(22, 8),
    to_signed(24, 8),
    to_signed(11, 8),
    to_signed(-15, 8),
    to_signed(-45, 8),
    to_signed(-67, 8),
    to_signed(-75, 8),
    to_signed(-70, 8),
    to_signed(-55, 8),
    to_signed(-33, 8),
    to_signed(-7, 8),
    to_signed(16, 8),
    to_signed(33, 8),
    to_signed(42, 8),
    to_signed(42, 8),
    to_signed(36, 8),
    to_signed(27, 8),
    to_signed(16, 8),
    to_signed(3, 8),
    to_signed(-9, 8),
    to_signed(-17, 8),
    to_signed(-21, 8),
    to_signed(-21, 8),
    to_signed(-18, 8),
    to_signed(-12, 8),
    to_signed(-3, 8),
    to_signed(7, 8),
    to_signed(17, 8),
    to_signed(23, 8),
    to_signed(23, 8),
    to_signed(16, 8),
    to_signed(0, 8),
    to_signed(-19, 8),
    to_signed(-37, 8),
    to_signed(-48, 8),
    to_signed(-52, 8),
    to_signed(-47, 8),
    to_signed(-35, 8),
    to_signed(-18, 8),
    to_signed(1, 8),
    to_signed(19, 8),
    to_signed(31, 8),
    to_signed(37, 8),
    to_signed(38, 8),
    to_signed(38, 8),
    to_signed(34, 8),
    to_signed(25, 8),
    to_signed(12, 8),
    to_signed(-1, 8),
    to_signed(-8, 8),
    to_signed(-11, 8),
    to_signed(-9, 8),
    to_signed(-5, 8),
    to_signed(3, 8),
    to_signed(15, 8),
    to_signed(29, 8),
    to_signed(41, 8),
    to_signed(47, 8),
    to_signed(49, 8),
    to_signed(47, 8),
    to_signed(42, 8),
    to_signed(31, 8),
    to_signed(13, 8),
    to_signed(-7, 8),
    to_signed(-30, 8),
    to_signed(-54, 8),
    to_signed(-78, 8),
    to_signed(-93, 8),
    to_signed(-94, 8),
    to_signed(-80, 8),
    to_signed(-54, 8),
    to_signed(-25, 8),
    to_signed(1, 8),
    to_signed(21, 8),
    to_signed(31, 8),
    to_signed(29, 8),
    to_signed(13, 8),
    to_signed(-13, 8),
    to_signed(-37, 8),
    to_signed(-51, 8),
    to_signed(-52, 8),
    to_signed(-44, 8),
    to_signed(-29, 8),
    to_signed(-8, 8),
    to_signed(16, 8),
    to_signed(37, 8),
    to_signed(52, 8),
    to_signed(58, 8),
    to_signed(57, 8),
    to_signed(50, 8),
    to_signed(39, 8),
    to_signed(24, 8),
    to_signed(9, 8),
    to_signed(-4, 8),
    to_signed(-11, 8),
    to_signed(-14, 8),
    to_signed(-14, 8),
    to_signed(-13, 8),
    to_signed(-7, 8),
    to_signed(2, 8),
    to_signed(12, 8),
    to_signed(19, 8),
    to_signed(22, 8),
    to_signed(16, 8),
    to_signed(4, 8),
    to_signed(-15, 8),
    to_signed(-33, 8),
    to_signed(-47, 8),
    to_signed(-53, 8),
    to_signed(-51, 8),
    to_signed(-41, 8),
    to_signed(-25, 8),
    to_signed(-6, 8),
    to_signed(14, 8),
    to_signed(29, 8),
    to_signed(38, 8),
    to_signed(42, 8),
    to_signed(42, 8),
    to_signed(41, 8),
    to_signed(35, 8),
    to_signed(24, 8),
    to_signed(11, 8),
    to_signed(3, 8),
    to_signed(-1, 8),
    to_signed(-1, 8),
    to_signed(0, 8),
    to_signed(5, 8),
    to_signed(15, 8),
    to_signed(30, 8),
    to_signed(45, 8),
    to_signed(55, 8),
    to_signed(59, 8),
    to_signed(58, 8),
    to_signed(54, 8),
    to_signed(46, 8),
    to_signed(31, 8),
    to_signed(11, 8),
    to_signed(-11, 8),
    to_signed(-33, 8),
    to_signed(-54, 8),
    to_signed(-73, 8),
    to_signed(-83, 8),
    to_signed(-80, 8),
    to_signed(-63, 8),
    to_signed(-38, 8),
    to_signed(-12, 8),
    to_signed(9, 8),
    to_signed(23, 8),
    to_signed(29, 8),
    to_signed(24, 8),
    to_signed(6, 8),
    to_signed(-17, 8),
    to_signed(-37, 8),
    to_signed(-48, 8),
    to_signed(-49, 8),
    to_signed(-41, 8),
    to_signed(-26, 8),
    to_signed(-5, 8),
    to_signed(18, 8),
    to_signed(38, 8),
    to_signed(51, 8),
    to_signed(55, 8),
    to_signed(50, 8),
    to_signed(39, 8),
    to_signed(25, 8),
    to_signed(9, 8),
    to_signed(-7, 8),
    to_signed(-18, 8),
    to_signed(-24, 8),
    to_signed(-25, 8),
    to_signed(-23, 8),
    to_signed(-16, 8),
    to_signed(-6, 8),
    to_signed(4, 8),
    to_signed(11, 8),
    to_signed(13, 8),
    to_signed(12, 8),
    to_signed(6, 8),
    to_signed(-7, 8),
    to_signed(-23, 8),
    to_signed(-39, 8),
    to_signed(-51, 8),
    to_signed(-55, 8),
    to_signed(-51, 8),
    to_signed(-40, 8),
    to_signed(-24, 8),
    to_signed(-5, 8),
    to_signed(13, 8),
    to_signed(29, 8),
    to_signed(37, 8),
    to_signed(39, 8),
    to_signed(38, 8),
    to_signed(35, 8),
    to_signed(29, 8),
    to_signed(18, 8),
    to_signed(6, 8),
    to_signed(-1, 8),
    to_signed(-3, 8),
    to_signed(-2, 8),
    to_signed(3, 8),
    to_signed(10, 8),
    to_signed(21, 8),
    to_signed(36, 8),
    to_signed(51, 8),
    to_signed(61, 8),
    to_signed(63, 8),
    to_signed(60, 8),
    to_signed(53, 8),
    to_signed(42, 8),
    to_signed(26, 8),
    to_signed(7, 8),
    to_signed(-15, 8),
    to_signed(-37, 8),
    to_signed(-60, 8),
    to_signed(-77, 8),
    to_signed(-83, 8),
    to_signed(-74, 8),
    to_signed(-53, 8),
    to_signed(-26, 8),
    to_signed(1, 8),
    to_signed(21, 8),
    to_signed(32, 8),
    to_signed(32, 8),
    to_signed(18, 8),
    to_signed(-5, 8),
    to_signed(-30, 8),
    to_signed(-49, 8),
    to_signed(-57, 8),
    to_signed(-55, 8),
    to_signed(-43, 8),
    to_signed(-22, 8),
    to_signed(3, 8),
    to_signed(28, 8),
    to_signed(45, 8),
    to_signed(53, 8),
    to_signed(53, 8),
    to_signed(47, 8),
    to_signed(38, 8),
    to_signed(26, 8),
    to_signed(11, 8),
    to_signed(-5, 8),
    to_signed(-19, 8),
    to_signed(-27, 8),
    to_signed(-31, 8),
    to_signed(-30, 8),
    to_signed(-22, 8),
    to_signed(-10, 8),
    to_signed(3, 8),
    to_signed(13, 8),
    to_signed(16, 8),
    to_signed(14, 8),
    to_signed(4, 8),
    to_signed(-13, 8),
    to_signed(-34, 8),
    to_signed(-54, 8),
    to_signed(-65, 8),
    to_signed(-66, 8),
    to_signed(-57, 8),
    to_signed(-41, 8),
    to_signed(-22, 8),
    to_signed(-2, 8),
    to_signed(15, 8),
    to_signed(27, 8),
    to_signed(32, 8),
    to_signed(34, 8),
    to_signed(34, 8),
    to_signed(32, 8),
    to_signed(25, 8),
    to_signed(14, 8),
    to_signed(4, 8),
    to_signed(-2, 8),
    to_signed(-3, 8),
    to_signed(0, 8),
    to_signed(5, 8),
    to_signed(14, 8),
    to_signed(27, 8),
    to_signed(43, 8),
    to_signed(57, 8),
    to_signed(64, 8),
    to_signed(64, 8),
    to_signed(60, 8),
    to_signed(52, 8),
    to_signed(39, 8),
    to_signed(21, 8),
    to_signed(1, 8),
    to_signed(-19, 8),
    to_signed(-40, 8),
    to_signed(-59, 8),
    to_signed(-74, 8),
    to_signed(-78, 8),
    to_signed(-69, 8),
    to_signed(-50, 8),
    to_signed(-25, 8),
    to_signed(-1, 8),
    to_signed(17, 8),
    to_signed(27, 8),
    to_signed(24, 8),
    to_signed(8, 8),
    to_signed(-18, 8),
    to_signed(-45, 8),
    to_signed(-63, 8),
    to_signed(-68, 8),
    to_signed(-62, 8),
    to_signed(-45, 8),
    to_signed(-23, 8),
    to_signed(1, 8),
    to_signed(21, 8),
    to_signed(34, 8),
    to_signed(38, 8),
    to_signed(36, 8),
    to_signed(30, 8),
    to_signed(23, 8),
    to_signed(13, 8),
    to_signed(0, 8),
    to_signed(-12, 8),
    to_signed(-23, 8),
    to_signed(-29, 8),
    to_signed(-32, 8),
    to_signed(-31, 8),
    to_signed(-23, 8),
    to_signed(-12, 8),
    to_signed(-2, 8),
    to_signed(6, 8),
    to_signed(9, 8),
    to_signed(7, 8),
    to_signed(-3, 8),
    to_signed(-19, 8),
    to_signed(-39, 8),
    to_signed(-55, 8),
    to_signed(-64, 8),
    to_signed(-63, 8),
    to_signed(-52, 8),
    to_signed(-36, 8),
    to_signed(-17, 8),
    to_signed(2, 8),
    to_signed(18, 8),
    to_signed(28, 8),
    to_signed(32, 8),
    to_signed(32, 8),
    to_signed(31, 8),
    to_signed(28, 8),
    to_signed(23, 8),
    to_signed(16, 8),
    to_signed(9, 8),
    to_signed(5, 8),
    to_signed(4, 8),
    to_signed(6, 8),
    to_signed(11, 8),
    to_signed(21, 8),
    to_signed(33, 8),
    to_signed(46, 8),
    to_signed(56, 8),
    to_signed(60, 8),
    to_signed(62, 8),
    to_signed(62, 8),
    to_signed(57, 8),
    to_signed(46, 8),
    to_signed(29, 8),
    to_signed(9, 8),
    to_signed(-12, 8),
    to_signed(-35, 8),
    to_signed(-57, 8),
    to_signed(-73, 8),
    to_signed(-76, 8),
    to_signed(-67, 8),
    to_signed(-46, 8),
    to_signed(-20, 8),
    to_signed(4, 8),
    to_signed(22, 8),
    to_signed(31, 8),
    to_signed(27, 8),
    to_signed(8, 8),
    to_signed(-19, 8),
    to_signed(-44, 8),
    to_signed(-58, 8),
    to_signed(-60, 8),
    to_signed(-51, 8),
    to_signed(-34, 8),
    to_signed(-12, 8),
    to_signed(11, 8),
    to_signed(30, 8),
    to_signed(42, 8),
    to_signed(46, 8),
    to_signed(44, 8),
    to_signed(36, 8),
    to_signed(27, 8),
    to_signed(16, 8),
    to_signed(3, 8),
    to_signed(-9, 8),
    to_signed(-17, 8),
    to_signed(-21, 8),
    to_signed(-22, 8),
    to_signed(-18, 8),
    to_signed(-10, 8),
    to_signed(1, 8),
    to_signed(11, 8),
    to_signed(19, 8),
    to_signed(22, 8),
    to_signed(18, 8),
    to_signed(6, 8),
    to_signed(-12, 8),
    to_signed(-29, 8),
    to_signed(-41, 8),
    to_signed(-46, 8),
    to_signed(-41, 8),
    to_signed(-29, 8),
    to_signed(-14, 8),
    to_signed(3, 8),
    to_signed(19, 8),
    to_signed(32, 8),
    to_signed(39, 8),
    to_signed(41, 8),
    to_signed(42, 8),
    to_signed(41, 8),
    to_signed(37, 8),
    to_signed(30, 8),
    to_signed(22, 8),
    to_signed(16, 8),
    to_signed(15, 8),
    to_signed(15, 8),
    to_signed(17, 8),
    to_signed(21, 8),
    to_signed(27, 8),
    to_signed(37, 8),
    to_signed(48, 8),
    to_signed(55, 8),
    to_signed(58, 8),
    to_signed(58, 8),
    to_signed(57, 8),
    to_signed(51, 8),
    to_signed(38, 8),
    to_signed(20, 8),
    to_signed(-1, 8),
    to_signed(-22, 8),
    to_signed(-45, 8),
    to_signed(-67, 8),
    to_signed(-82, 8),
    to_signed(-84, 8),
    to_signed(-71, 8),
    to_signed(-47, 8),
    to_signed(-19, 8),
    to_signed(5, 8),
    to_signed(22, 8),
    to_signed(28, 8),
    to_signed(23, 8),
    to_signed(4, 8),
    to_signed(-21, 8),
    to_signed(-44, 8),
    to_signed(-56, 8),
    to_signed(-57, 8),
    to_signed(-49, 8),
    to_signed(-32, 8),
    to_signed(-10, 8),
    to_signed(13, 8),
    to_signed(31, 8),
    to_signed(42, 8),
    to_signed(45, 8),
    to_signed(41, 8),
    to_signed(35, 8),
    to_signed(26, 8),
    to_signed(15, 8),
    to_signed(2, 8),
    to_signed(-10, 8),
    to_signed(-17, 8),
    to_signed(-22, 8),
    to_signed(-24, 8),
    to_signed(-21, 8),
    to_signed(-12, 8),
    to_signed(0, 8),
    to_signed(12, 8),
    to_signed(21, 8),
    to_signed(23, 8),
    to_signed(18, 8),
    to_signed(4, 8),
    to_signed(-16, 8),
    to_signed(-36, 8),
    to_signed(-50, 8),
    to_signed(-53, 8),
    to_signed(-44, 8),
    to_signed(-28, 8),
    to_signed(-10, 8),
    to_signed(7, 8),
    to_signed(22, 8),
    to_signed(34, 8),
    to_signed(40, 8),
    to_signed(41, 8),
    to_signed(39, 8),
    to_signed(35, 8),
    to_signed(27, 8),
    to_signed(16, 8),
    to_signed(7, 8),
    to_signed(1, 8),
    to_signed(-2, 8),
    to_signed(-2, 8),
    to_signed(-1, 8),
    to_signed(3, 8),
    to_signed(13, 8),
    to_signed(29, 8),
    to_signed(45, 8),
    to_signed(55, 8),
    to_signed(57, 8),
    to_signed(54, 8),
    to_signed(48, 8),
    to_signed(37, 8),
    to_signed(20, 8),
    to_signed(1, 8),
    to_signed(-16, 8),
    to_signed(-32, 8),
    to_signed(-50, 8),
    to_signed(-67, 8),
    to_signed(-80, 8),
    to_signed(-81, 8),
    to_signed(-68, 8),
    to_signed(-45, 8),
    to_signed(-19, 8),
    to_signed(2, 8),
    to_signed(16, 8),
    to_signed(22, 8),
    to_signed(17, 8),
    to_signed(-1, 8),
    to_signed(-26, 8),
    to_signed(-48, 8),
    to_signed(-59, 8),
    to_signed(-60, 8),
    to_signed(-52, 8),
    to_signed(-36, 8),
    to_signed(-13, 8),
    to_signed(11, 8),
    to_signed(30, 8),
    to_signed(41, 8),
    to_signed(41, 8),
    to_signed(35, 8),
    to_signed(27, 8),
    to_signed(17, 8),
    to_signed(5, 8),
    to_signed(-9, 8),
    to_signed(-19, 8),
    to_signed(-23, 8),
    to_signed(-24, 8),
    to_signed(-24, 8),
    to_signed(-22, 8),
    to_signed(-16, 8),
    to_signed(-7, 8),
    to_signed(3, 8),
    to_signed(12, 8),
    to_signed(15, 8),
    to_signed(12, 8),
    to_signed(0, 8),
    to_signed(-19, 8),
    to_signed(-38, 8),
    to_signed(-53, 8),
    to_signed(-57, 8),
    to_signed(-49, 8),
    to_signed(-35, 8),
    to_signed(-20, 8),
    to_signed(-3, 8),
    to_signed(13, 8),
    to_signed(26, 8),
    to_signed(32, 8),
    to_signed(33, 8),
    to_signed(32, 8),
    to_signed(28, 8),
    to_signed(23, 8),
    to_signed(16, 8),
    to_signed(10, 8),
    to_signed(5, 8),
    to_signed(2, 8),
    to_signed(1, 8),
    to_signed(2, 8),
    to_signed(6, 8),
    to_signed(16, 8),
    to_signed(32, 8),
    to_signed(48, 8),
    to_signed(59, 8),
    to_signed(63, 8),
    to_signed(64, 8),
    to_signed(62, 8),
    to_signed(52, 8),
    to_signed(34, 8),
    to_signed(12, 8),
    to_signed(-8, 8),
    to_signed(-27, 8),
    to_signed(-46, 8),
    to_signed(-66, 8),
    to_signed(-81, 8),
    to_signed(-83, 8),
    to_signed(-69, 8),
    to_signed(-44, 8),
    to_signed(-17, 8),
    to_signed(3, 8),
    to_signed(16, 8),
    to_signed(22, 8),
    to_signed(17, 8),
    to_signed(0, 8),
    to_signed(-25, 8),
    to_signed(-48, 8),
    to_signed(-60, 8),
    to_signed(-62, 8),
    to_signed(-53, 8),
    to_signed(-38, 8),
    to_signed(-18, 8),
    to_signed(3, 8),
    to_signed(21, 8),
    to_signed(31, 8),
    to_signed(33, 8),
    to_signed(30, 8),
    to_signed(25, 8),
    to_signed(17, 8),
    to_signed(5, 8),
    to_signed(-8, 8),
    to_signed(-19, 8),
    to_signed(-26, 8),
    to_signed(-31, 8),
    to_signed(-33, 8),
    to_signed(-32, 8),
    to_signed(-25, 8),
    to_signed(-13, 8),
    to_signed(0, 8),
    to_signed(10, 8),
    to_signed(13, 8),
    to_signed(10, 8),
    to_signed(-1, 8),
    to_signed(-16, 8),
    to_signed(-33, 8),
    to_signed(-45, 8),
    to_signed(-48, 8),
    to_signed(-42, 8),
    to_signed(-29, 8),
    to_signed(-14, 8),
    to_signed(4, 8),
    to_signed(21, 8),
    to_signed(34, 8),
    to_signed(40, 8),
    to_signed(39, 8),
    to_signed(36, 8),
    to_signed(32, 8),
    to_signed(27, 8),
    to_signed(22, 8),
    to_signed(15, 8),
    to_signed(10, 8),
    to_signed(7, 8),
    to_signed(6, 8),
    to_signed(7, 8),
    to_signed(12, 8),
    to_signed(21, 8),
    to_signed(34, 8),
    to_signed(47, 8),
    to_signed(55, 8),
    to_signed(59, 8),
    to_signed(60, 8),
    to_signed(59, 8),
    to_signed(51, 8),
    to_signed(35, 8),
    to_signed(14, 8),
    to_signed(-7, 8),
    to_signed(-28, 8),
    to_signed(-50, 8),
    to_signed(-72, 8),
    to_signed(-86, 8),
    to_signed(-85, 8),
    to_signed(-65, 8),
    to_signed(-36, 8),
    to_signed(-9, 8),
    to_signed(10, 8),
    to_signed(22, 8),
    to_signed(25, 8),
    to_signed(17, 8),
    to_signed(-5, 8),
    to_signed(-33, 8),
    to_signed(-56, 8),
    to_signed(-66, 8),
    to_signed(-61, 8),
    to_signed(-47, 8),
    to_signed(-29, 8),
    to_signed(-10, 8),
    to_signed(10, 8),
    to_signed(26, 8),
    to_signed(34, 8),
    to_signed(33, 8),
    to_signed(28, 8),
    to_signed(22, 8),
    to_signed(14, 8),
    to_signed(5, 8),
    to_signed(-6, 8),
    to_signed(-15, 8),
    to_signed(-21, 8),
    to_signed(-24, 8),
    to_signed(-24, 8),
    to_signed(-20, 8),
    to_signed(-12, 8),
    to_signed(0, 8),
    to_signed(13, 8),
    to_signed(21, 8),
    to_signed(23, 8),
    to_signed(18, 8),
    to_signed(6, 8),
    to_signed(-9, 8),
    to_signed(-24, 8),
    to_signed(-34, 8),
    to_signed(-35, 8),
    to_signed(-28, 8),
    to_signed(-16, 8),
    to_signed(-1, 8),
    to_signed(16, 8),
    to_signed(34, 8),
    to_signed(46, 8),
    to_signed(51, 8),
    to_signed(49, 8),
    to_signed(46, 8),
    to_signed(42, 8),
    to_signed(36, 8),
    to_signed(26, 8),
    to_signed(15, 8),
    to_signed(8, 8),
    to_signed(4, 8),
    to_signed(5, 8),
    to_signed(8, 8),
    to_signed(14, 8),
    to_signed(24, 8),
    to_signed(38, 8),
    to_signed(49, 8),
    to_signed(55, 8),
    to_signed(56, 8),
    to_signed(55, 8),
    to_signed(53, 8),
    to_signed(46, 8),
    to_signed(32, 8),
    to_signed(12, 8),
    to_signed(-9, 8),
    to_signed(-31, 8),
    to_signed(-55, 8),
    to_signed(-75, 8),
    to_signed(-86, 8),
    to_signed(-81, 8),
    to_signed(-61, 8),
    to_signed(-34, 8),
    to_signed(-10, 8),
    to_signed(6, 8),
    to_signed(15, 8),
    to_signed(17, 8),
    to_signed(9, 8),
    to_signed(-11, 8),
    to_signed(-35, 8),
    to_signed(-53, 8),
    to_signed(-57, 8),
    to_signed(-50, 8),
    to_signed(-37, 8),
    to_signed(-19, 8),
    to_signed(1, 8),
    to_signed(20, 8),
    to_signed(33, 8),
    to_signed(39, 8),
    to_signed(37, 8),
    to_signed(30, 8),
    to_signed(23, 8),
    to_signed(16, 8),
    to_signed(7, 8),
    to_signed(-2, 8),
    to_signed(-9, 8),
    to_signed(-14, 8),
    to_signed(-16, 8),
    to_signed(-17, 8),
    to_signed(-14, 8),
    to_signed(-6, 8),
    to_signed(4, 8),
    to_signed(12, 8),
    to_signed(17, 8),
    to_signed(15, 8),
    to_signed(9, 8),
    to_signed(-3, 8),
    to_signed(-17, 8),
    to_signed(-29, 8),
    to_signed(-36, 8),
    to_signed(-36, 8),
    to_signed(-28, 8),
    to_signed(-16, 8),
    to_signed(-2, 8),
    to_signed(13, 8),
    to_signed(27, 8),
    to_signed(36, 8),
    to_signed(38, 8),
    to_signed(36, 8),
    to_signed(33, 8),
    to_signed(30, 8),
    to_signed(24, 8),
    to_signed(17, 8),
    to_signed(10, 8),
    to_signed(7, 8),
    to_signed(6, 8),
    to_signed(8, 8),
    to_signed(11, 8),
    to_signed(17, 8),
    to_signed(27, 8),
    to_signed(41, 8),
    to_signed(52, 8),
    to_signed(58, 8),
    to_signed(59, 8),
    to_signed(59, 8),
    to_signed(55, 8),
    to_signed(44, 8),
    to_signed(25, 8),
    to_signed(3, 8),
    to_signed(-19, 8),
    to_signed(-41, 8),
    to_signed(-63, 8),
    to_signed(-81, 8),
    to_signed(-86, 8),
    to_signed(-75, 8),
    to_signed(-50, 8),
    to_signed(-22, 8),
    to_signed(0, 8),
    to_signed(12, 8),
    to_signed(16, 8),
    to_signed(12, 8),
    to_signed(-4, 8),
    to_signed(-28, 8),
    to_signed(-51, 8),
    to_signed(-62, 8),
    to_signed(-60, 8),
    to_signed(-48, 8),
    to_signed(-32, 8),
    to_signed(-13, 8),
    to_signed(8, 8),
    to_signed(26, 8),
    to_signed(37, 8),
    to_signed(40, 8),
    to_signed(35, 8),
    to_signed(26, 8),
    to_signed(17, 8),
    to_signed(6, 8),
    to_signed(-8, 8),
    to_signed(-21, 8),
    to_signed(-29, 8),
    to_signed(-32, 8),
    to_signed(-32, 8),
    to_signed(-29, 8),
    to_signed(-22, 8),
    to_signed(-12, 8),
    to_signed(-2, 8),
    to_signed(4, 8),
    to_signed(7, 8),
    to_signed(4, 8),
    to_signed(-2, 8),
    to_signed(-13, 8),
    to_signed(-26, 8),
    to_signed(-38, 8),
    to_signed(-44, 8),
    to_signed(-42, 8),
    to_signed(-33, 8),
    to_signed(-20, 8),
    to_signed(-5, 8),
    to_signed(11, 8),
    to_signed(27, 8),
    to_signed(36, 8),
    to_signed(38, 8),
    to_signed(35, 8),
    to_signed(32, 8),
    to_signed(28, 8),
    to_signed(22, 8),
    to_signed(14, 8),
    to_signed(9, 8),
    to_signed(6, 8),
    to_signed(6, 8),
    to_signed(7, 8),
    to_signed(10, 8),
    to_signed(16, 8),
    to_signed(28, 8),
    to_signed(42, 8),
    to_signed(52, 8),
    to_signed(55, 8),
    to_signed(54, 8),
    to_signed(52, 8),
    to_signed(46, 8),
    to_signed(33, 8),
    to_signed(15, 8),
    to_signed(-5, 8),
    to_signed(-23, 8),
    to_signed(-42, 8),
    to_signed(-62, 8),
    to_signed(-78, 8),
    to_signed(-80, 8),
    to_signed(-67, 8),
    to_signed(-42, 8),
    to_signed(-17, 8),
    to_signed(1, 8),
    to_signed(10, 8),
    to_signed(13, 8),
    to_signed(8, 8),
    to_signed(-9, 8),
    to_signed(-32, 8),
    to_signed(-50, 8),
    to_signed(-55, 8),
    to_signed(-47, 8),
    to_signed(-33, 8),
    to_signed(-16, 8),
    to_signed(1, 8),
    to_signed(17, 8),
    to_signed(31, 8),
    to_signed(37, 8),
    to_signed(36, 8),
    to_signed(28, 8),
    to_signed(20, 8),
    to_signed(11, 8),
    to_signed(0, 8),
    to_signed(-13, 8),
    to_signed(-23, 8),
    to_signed(-28, 8),
    to_signed(-29, 8),
    to_signed(-28, 8),
    to_signed(-26, 8),
    to_signed(-21, 8),
    to_signed(-14, 8),
    to_signed(-7, 8),
    to_signed(-2, 8),
    to_signed(1, 8),
    to_signed(0, 8),
    to_signed(-6, 8),
    to_signed(-16, 8),
    to_signed(-27, 8),
    to_signed(-36, 8),
    to_signed(-37, 8),
    to_signed(-30, 8),
    to_signed(-19, 8),
    to_signed(-8, 8),
    to_signed(3, 8),
    to_signed(16, 8),
    to_signed(28, 8),
    to_signed(35, 8),
    to_signed(35, 8),
    to_signed(33, 8),
    to_signed(30, 8),
    to_signed(28, 8),
    to_signed(24, 8),
    to_signed(17, 8),
    to_signed(12, 8),
    to_signed(8, 8),
    to_signed(8, 8),
    to_signed(9, 8),
    to_signed(12, 8),
    to_signed(18, 8),
    to_signed(29, 8),
    to_signed(43, 8),
    to_signed(53, 8),
    to_signed(58, 8),
    to_signed(59, 8),
    to_signed(57, 8),
    to_signed(50, 8),
    to_signed(36, 8),
    to_signed(17, 8),
    to_signed(-3, 8),
    to_signed(-23, 8),
    to_signed(-44, 8),
    to_signed(-65, 8),
    to_signed(-77, 8),
    to_signed(-74, 8),
    to_signed(-56, 8),
    to_signed(-31, 8),
    to_signed(-9, 8),
    to_signed(7, 8),
    to_signed(16, 8),
    to_signed(19, 8),
    to_signed(12, 8),
    to_signed(-8, 8),
    to_signed(-35, 8),
    to_signed(-54, 8),
    to_signed(-58, 8),
    to_signed(-51, 8),
    to_signed(-37, 8),
    to_signed(-20, 8),
    to_signed(1, 8),
    to_signed(21, 8),
    to_signed(36, 8),
    to_signed(41, 8),
    to_signed(36, 8),
    to_signed(26, 8),
    to_signed(17, 8),
    to_signed(7, 8),
    to_signed(-4, 8),
    to_signed(-16, 8),
    to_signed(-23, 8),
    to_signed(-25, 8),
    to_signed(-23, 8),
    to_signed(-22, 8),
    to_signed(-20, 8),
    to_signed(-14, 8),
    to_signed(-5, 8),
    to_signed(5, 8),
    to_signed(13, 8),
    to_signed(18, 8),
    to_signed(18, 8),
    to_signed(10, 8),
    to_signed(-3, 8),
    to_signed(-18, 8),
    to_signed(-29, 8),
    to_signed(-31, 8),
    to_signed(-25, 8),
    to_signed(-14, 8),
    to_signed(0, 8),
    to_signed(15, 8),
    to_signed(31, 8),
    to_signed(43, 8),
    to_signed(47, 8),
    to_signed(45, 8),
    to_signed(41, 8),
    to_signed(37, 8),
    to_signed(33, 8),
    to_signed(27, 8),
    to_signed(20, 8),
    to_signed(16, 8),
    to_signed(15, 8),
    to_signed(17, 8),
    to_signed(19, 8),
    to_signed(22, 8),
    to_signed(28, 8),
    to_signed(38, 8),
    to_signed(48, 8),
    to_signed(55, 8),
    to_signed(58, 8),
    to_signed(59, 8),
    to_signed(57, 8),
    to_signed(51, 8),
    to_signed(37, 8),
    to_signed(18, 8),
    to_signed(-3, 8),
    to_signed(-25, 8),
    to_signed(-50, 8),
    to_signed(-73, 8),
    to_signed(-84, 8),
    to_signed(-78, 8),
    to_signed(-57, 8),
    to_signed(-30, 8),
    to_signed(-6, 8),
    to_signed(10, 8),
    to_signed(19, 8),
    to_signed(20, 8),
    to_signed(7, 8),
    to_signed(-17, 8),
    to_signed(-44, 8),
    to_signed(-61, 8),
    to_signed(-65, 8),
    to_signed(-58, 8),
    to_signed(-45, 8),
    to_signed(-27, 8),
    to_signed(-3, 8),
    to_signed(21, 8),
    to_signed(37, 8),
    to_signed(42, 8),
    to_signed(36, 8),
    to_signed(26, 8),
    to_signed(16, 8),
    to_signed(4, 8),
    to_signed(-10, 8),
    to_signed(-22, 8),
    to_signed(-29, 8),
    to_signed(-29, 8),
    to_signed(-28, 8),
    to_signed(-25, 8),
    to_signed(-21, 8),
    to_signed(-13, 8),
    to_signed(-3, 8),
    to_signed(7, 8),
    to_signed(13, 8),
    to_signed(15, 8),
    to_signed(13, 8),
    to_signed(4, 8),
    to_signed(-9, 8),
    to_signed(-24, 8),
    to_signed(-32, 8),
    to_signed(-32, 8),
    to_signed(-24, 8),
    to_signed(-13, 8),
    to_signed(-1, 8),
    to_signed(12, 8),
    to_signed(26, 8),
    to_signed(37, 8),
    to_signed(41, 8),
    to_signed(40, 8),
    to_signed(38, 8),
    to_signed(35, 8),
    to_signed(28, 8),
    to_signed(20, 8),
    to_signed(10, 8),
    to_signed(4, 8),
    to_signed(2, 8),
    to_signed(4, 8),
    to_signed(7, 8),
    to_signed(14, 8),
    to_signed(25, 8),
    to_signed(38, 8),
    to_signed(49, 8),
    to_signed(54, 8),
    to_signed(56, 8),
    to_signed(56, 8),
    to_signed(52, 8),
    to_signed(42, 8),
    to_signed(26, 8),
    to_signed(8, 8),
    to_signed(-12, 8),
    to_signed(-36, 8),
    to_signed(-62, 8),
    to_signed(-83, 8),
    to_signed(-88, 8),
    to_signed(-74, 8),
    to_signed(-47, 8),
    to_signed(-18, 8),
    to_signed(3, 8),
    to_signed(16, 8),
    to_signed(20, 8),
    to_signed(14, 8),
    to_signed(-6, 8),
    to_signed(-34, 8),
    to_signed(-58, 8),
    to_signed(-69, 8),
    to_signed(-66, 8),
    to_signed(-55, 8),
    to_signed(-39, 8),
    to_signed(-17, 8),
    to_signed(8, 8),
    to_signed(29, 8),
    to_signed(40, 8),
    to_signed(40, 8),
    to_signed(31, 8),
    to_signed(19, 8),
    to_signed(6, 8),
    to_signed(-9, 8),
    to_signed(-23, 8),
    to_signed(-34, 8),
    to_signed(-36, 8),
    to_signed(-35, 8),
    to_signed(-32, 8),
    to_signed(-29, 8),
    to_signed(-23, 8),
    to_signed(-14, 8),
    to_signed(-4, 8),
    to_signed(4, 8),
    to_signed(10, 8),
    to_signed(11, 8),
    to_signed(6, 8),
    to_signed(-5, 8),
    to_signed(-21, 8),
    to_signed(-35, 8),
    to_signed(-41, 8),
    to_signed(-37, 8),
    to_signed(-27, 8),
    to_signed(-16, 8),
    to_signed(-4, 8),
    to_signed(10, 8),
    to_signed(23, 8),
    to_signed(32, 8),
    to_signed(34, 8),
    to_signed(33, 8),
    to_signed(30, 8),
    to_signed(27, 8),
    to_signed(22, 8),
    to_signed(16, 8),
    to_signed(9, 8),
    to_signed(4, 8),
    to_signed(3, 8),
    to_signed(4, 8),
    to_signed(9, 8),
    to_signed(17, 8),
    to_signed(31, 8),
    to_signed(46, 8),
    to_signed(58, 8),
    to_signed(65, 8),
    to_signed(69, 8),
    to_signed(69, 8),
    to_signed(62, 8),
    to_signed(47, 8),
    to_signed(27, 8),
    to_signed(4, 8),
    to_signed(-22, 8),
    to_signed(-50, 8),
    to_signed(-76, 8),
    to_signed(-89, 8),
    to_signed(-85, 8),
    to_signed(-63, 8),
    to_signed(-33, 8),
    to_signed(-6, 8),
    to_signed(12, 8),
    to_signed(21, 8),
    to_signed(19, 8),
    to_signed(4, 8),
    to_signed(-24, 8),
    to_signed(-54, 8),
    to_signed(-73, 8),
    to_signed(-79, 8),
    to_signed(-72, 8),
    to_signed(-59, 8),
    to_signed(-40, 8),
    to_signed(-17, 8),
    to_signed(6, 8),
    to_signed(25, 8),
    to_signed(33, 8),
    to_signed(31, 8),
    to_signed(23, 8),
    to_signed(12, 8),
    to_signed(-1, 8),
    to_signed(-18, 8),
    to_signed(-33, 8),
    to_signed(-42, 8),
    to_signed(-42, 8),
    to_signed(-39, 8),
    to_signed(-35, 8),
    to_signed(-30, 8),
    to_signed(-20, 8),
    to_signed(-8, 8),
    to_signed(4, 8),
    to_signed(13, 8),
    to_signed(17, 8),
    to_signed(16, 8),
    to_signed(8, 8),
    to_signed(-5, 8),
    to_signed(-22, 8),
    to_signed(-36, 8),
    to_signed(-40, 8),
    to_signed(-34, 8),
    to_signed(-21, 8),
    to_signed(-6, 8),
    to_signed(10, 8),
    to_signed(27, 8),
    to_signed(41, 8),
    to_signed(49, 8),
    to_signed(51, 8),
    to_signed(48, 8),
    to_signed(42, 8),
    to_signed(34, 8),
    to_signed(26, 8),
    to_signed(18, 8),
    to_signed(13, 8),
    to_signed(10, 8),
    to_signed(11, 8),
    to_signed(16, 8),
    to_signed(24, 8),
    to_signed(35, 8),
    to_signed(48, 8),
    to_signed(59, 8),
    to_signed(67, 8),
    to_signed(71, 8),
    to_signed(72, 8),
    to_signed(67, 8),
    to_signed(54, 8),
    to_signed(34, 8),
    to_signed(12, 8),
    to_signed(-12, 8),
    to_signed(-37, 8),
    to_signed(-62, 8),
    to_signed(-81, 8),
    to_signed(-85, 8),
    to_signed(-72, 8),
    to_signed(-47, 8),
    to_signed(-20, 8),
    to_signed(-1, 8),
    to_signed(9, 8),
    to_signed(10, 8),
    to_signed(2, 8),
    to_signed(-18, 8),
    to_signed(-44, 8),
    to_signed(-67, 8),
    to_signed(-77, 8),
    to_signed(-74, 8),
    to_signed(-61, 8),
    to_signed(-43, 8),
    to_signed(-22, 8),
    to_signed(1, 8),
    to_signed(20, 8),
    to_signed(32, 8),
    to_signed(32, 8),
    to_signed(24, 8),
    to_signed(14, 8),
    to_signed(4, 8),
    to_signed(-6, 8),
    to_signed(-17, 8),
    to_signed(-25, 8),
    to_signed(-28, 8),
    to_signed(-27, 8),
    to_signed(-26, 8),
    to_signed(-24, 8),
    to_signed(-19, 8),
    to_signed(-12, 8),
    to_signed(-3, 8),
    to_signed(5, 8),
    to_signed(11, 8),
    to_signed(14, 8),
    to_signed(11, 8),
    to_signed(3, 8),
    to_signed(-8, 8),
    to_signed(-19, 8),
    to_signed(-25, 8),
    to_signed(-24, 8),
    to_signed(-16, 8),
    to_signed(-5, 8),
    to_signed(6, 8),
    to_signed(19, 8),
    to_signed(31, 8),
    to_signed(41, 8),
    to_signed(47, 8),
    to_signed(51, 8),
    to_signed(52, 8),
    to_signed(49, 8),
    to_signed(41, 8),
    to_signed(31, 8),
    to_signed(22, 8),
    to_signed(14, 8),
    to_signed(8, 8),
    to_signed(6, 8),
    to_signed(8, 8),
    to_signed(14, 8),
    to_signed(25, 8),
    to_signed(38, 8),
    to_signed(50, 8),
    to_signed(59, 8),
    to_signed(65, 8),
    to_signed(67, 8),
    to_signed(60, 8),
    to_signed(45, 8),
    to_signed(23, 8),
    to_signed(-1, 8),
    to_signed(-26, 8),
    to_signed(-53, 8),
    to_signed(-79, 8),
    to_signed(-94, 8),
    to_signed(-93, 8),
    to_signed(-74, 8),
    to_signed(-45, 8),
    to_signed(-19, 8),
    to_signed(-1, 8),
    to_signed(8, 8),
    to_signed(8, 8),
    to_signed(-3, 8),
    to_signed(-24, 8),
    to_signed(-49, 8),
    to_signed(-68, 8),
    to_signed(-73, 8),
    to_signed(-67, 8),
    to_signed(-54, 8),
    to_signed(-35, 8),
    to_signed(-13, 8),
    to_signed(9, 8),
    to_signed(28, 8),
    to_signed(39, 8),
    to_signed(40, 8),
    to_signed(34, 8),
    to_signed(26, 8),
    to_signed(17, 8),
    to_signed(5, 8),
    to_signed(-8, 8),
    to_signed(-18, 8),
    to_signed(-23, 8),
    to_signed(-23, 8),
    to_signed(-22, 8),
    to_signed(-17, 8),
    to_signed(-9, 8),
    to_signed(2, 8),
    to_signed(12, 8),
    to_signed(20, 8),
    to_signed(24, 8),
    to_signed(23, 8),
    to_signed(15, 8),
    to_signed(3, 8),
    to_signed(-11, 8),
    to_signed(-22, 8),
    to_signed(-27, 8),
    to_signed(-24, 8),
    to_signed(-15, 8),
    to_signed(-5, 8),
    to_signed(6, 8),
    to_signed(18, 8),
    to_signed(29, 8),
    to_signed(35, 8),
    to_signed(39, 8),
    to_signed(40, 8),
    to_signed(37, 8),
    to_signed(30, 8),
    to_signed(21, 8),
    to_signed(12, 8),
    to_signed(7, 8),
    to_signed(4, 8),
    to_signed(3, 8),
    to_signed(4, 8),
    to_signed(7, 8),
    to_signed(16, 8),
    to_signed(28, 8),
    to_signed(40, 8),
    to_signed(50, 8),
    to_signed(56, 8),
    to_signed(61, 8),
    to_signed(62, 8),
    to_signed(55, 8),
    to_signed(39, 8),
    to_signed(18, 8),
    to_signed(-4, 8),
    to_signed(-31, 8),
    to_signed(-60, 8),
    to_signed(-85, 8),
    to_signed(-97, 8),
    to_signed(-89, 8),
    to_signed(-64, 8),
    to_signed(-33, 8),
    to_signed(-7, 8),
    to_signed(9, 8),
    to_signed(15, 8),
    to_signed(12, 8),
    to_signed(-4, 8),
    to_signed(-29, 8),
    to_signed(-54, 8),
    to_signed(-69, 8),
    to_signed(-69, 8),
    to_signed(-59, 8),
    to_signed(-44, 8),
    to_signed(-25, 8),
    to_signed(-5, 8),
    to_signed(15, 8),
    to_signed(30, 8),
    to_signed(37, 8),
    to_signed(35, 8),
    to_signed(28, 8),
    to_signed(21, 8),
    to_signed(12, 8),
    to_signed(2, 8),
    to_signed(-9, 8),
    to_signed(-18, 8),
    to_signed(-23, 8),
    to_signed(-26, 8),
    to_signed(-26, 8),
    to_signed(-23, 8),
    to_signed(-16, 8),
    to_signed(-7, 8),
    to_signed(4, 8),
    to_signed(13, 8),
    to_signed(17, 8),
    to_signed(14, 8),
    to_signed(3, 8),
    to_signed(-11, 8),
    to_signed(-24, 8),
    to_signed(-33, 8),
    to_signed(-35, 8),
    to_signed(-30, 8),
    to_signed(-23, 8),
    to_signed(-14, 8),
    to_signed(-2, 8),
    to_signed(11, 8),
    to_signed(22, 8),
    to_signed(31, 8),
    to_signed(39, 8),
    to_signed(43, 8),
    to_signed(42, 8),
    to_signed(36, 8),
    to_signed(26, 8),
    to_signed(17, 8),
    to_signed(9, 8),
    to_signed(4, 8),
    to_signed(1, 8),
    to_signed(1, 8),
    to_signed(5, 8),
    to_signed(16, 8),
    to_signed(31, 8),
    to_signed(47, 8),
    to_signed(59, 8),
    to_signed(66, 8),
    to_signed(68, 8),
    to_signed(63, 8),
    to_signed(48, 8),
    to_signed(27, 8),
    to_signed(4, 8),
    to_signed(-20, 8),
    to_signed(-47, 8),
    to_signed(-72, 8),
    to_signed(-88, 8),
    to_signed(-89, 8),
    to_signed(-73, 8),
    to_signed(-44, 8),
    to_signed(-15, 8),
    to_signed(6, 8),
    to_signed(17, 8),
    to_signed(18, 8),
    to_signed(9, 8),
    to_signed(-11, 8),
    to_signed(-37, 8),
    to_signed(-59, 8),
    to_signed(-69, 8),
    to_signed(-66, 8),
    to_signed(-55, 8),
    to_signed(-37, 8),
    to_signed(-15, 8),
    to_signed(9, 8),
    to_signed(30, 8),
    to_signed(45, 8),
    to_signed(49, 8),
    to_signed(43, 8),
    to_signed(31, 8),
    to_signed(18, 8),
    to_signed(4, 8),
    to_signed(-10, 8),
    to_signed(-23, 8),
    to_signed(-30, 8),
    to_signed(-31, 8),
    to_signed(-29, 8),
    to_signed(-24, 8),
    to_signed(-17, 8),
    to_signed(-10, 8),
    to_signed(-1, 8),
    to_signed(8, 8),
    to_signed(14, 8),
    to_signed(14, 8),
    to_signed(6, 8),
    to_signed(-5, 8),
    to_signed(-16, 8),
    to_signed(-25, 8),
    to_signed(-28, 8),
    to_signed(-27, 8),
    to_signed(-21, 8),
    to_signed(-13, 8),
    to_signed(-3, 8),
    to_signed(9, 8),
    to_signed(20, 8),
    to_signed(30, 8),
    to_signed(38, 8),
    to_signed(44, 8),
    to_signed(47, 8),
    to_signed(44, 8),
    to_signed(36, 8),
    to_signed(27, 8),
    to_signed(18, 8),
    to_signed(10, 8),
    to_signed(4, 8),
    to_signed(0, 8),
    to_signed(0, 8),
    to_signed(7, 8),
    to_signed(21, 8),
    to_signed(39, 8),
    to_signed(56, 8),
    to_signed(69, 8),
    to_signed(76, 8),
    to_signed(74, 8),
    to_signed(63, 8),
    to_signed(43, 8),
    to_signed(18, 8),
    to_signed(-10, 8),
    to_signed(-39, 8),
    to_signed(-68, 8),
    to_signed(-90, 8),
    to_signed(-98, 8),
    to_signed(-88, 8),
    to_signed(-64, 8),
    to_signed(-34, 8),
    to_signed(-7, 8),
    to_signed(11, 8),
    to_signed(18, 8),
    to_signed(15, 8),
    to_signed(0, 8),
    to_signed(-23, 8),
    to_signed(-47, 8),
    to_signed(-63, 8),
    to_signed(-66, 8),
    to_signed(-59, 8),
    to_signed(-44, 8),
    to_signed(-24, 8),
    to_signed(0, 8),
    to_signed(24, 8),
    to_signed(45, 8),
    to_signed(56, 8),
    to_signed(56, 8),
    to_signed(48, 8),
    to_signed(36, 8),
    to_signed(23, 8),
    to_signed(8, 8),
    to_signed(-8, 8),
    to_signed(-23, 8),
    to_signed(-31, 8),
    to_signed(-33, 8),
    to_signed(-30, 8),
    to_signed(-23, 8),
    to_signed(-14, 8),
    to_signed(-3, 8),
    to_signed(10, 8),
    to_signed(22, 8),
    to_signed(27, 8),
    to_signed(22, 8),
    to_signed(10, 8),
    to_signed(-4, 8),
    to_signed(-16, 8),
    to_signed(-25, 8),
    to_signed(-29, 8),
    to_signed(-27, 8),
    to_signed(-20, 8),
    to_signed(-8, 8),
    to_signed(6, 8),
    to_signed(20, 8),
    to_signed(32, 8),
    to_signed(40, 8),
    to_signed(46, 8),
    to_signed(49, 8),
    to_signed(46, 8),
    to_signed(39, 8),
    to_signed(30, 8),
    to_signed(22, 8),
    to_signed(15, 8),
    to_signed(9, 8),
    to_signed(6, 8),
    to_signed(6, 8),
    to_signed(12, 8),
    to_signed(24, 8),
    to_signed(39, 8),
    to_signed(54, 8),
    to_signed(65, 8),
    to_signed(71, 8),
    to_signed(70, 8),
    to_signed(62, 8),
    to_signed(46, 8),
    to_signed(26, 8),
    to_signed(3, 8),
    to_signed(-24, 8),
    to_signed(-54, 8),
    to_signed(-80, 8),
    to_signed(-94, 8),
    to_signed(-91, 8),
    to_signed(-71, 8),
    to_signed(-41, 8),
    to_signed(-12, 8),
    to_signed(9, 8),
    to_signed(19, 8),
    to_signed(19, 8),
    to_signed(7, 8),
    to_signed(-15, 8),
    to_signed(-39, 8),
    to_signed(-56, 8),
    to_signed(-61, 8),
    to_signed(-55, 8),
    to_signed(-41, 8),
    to_signed(-23, 8),
    to_signed(-2, 8),
    to_signed(21, 8),
    to_signed(41, 8),
    to_signed(53, 8),
    to_signed(52, 8),
    to_signed(41, 8),
    to_signed(26, 8),
    to_signed(13, 8),
    to_signed(1, 8),
    to_signed(-11, 8),
    to_signed(-20, 8),
    to_signed(-26, 8),
    to_signed(-26, 8),
    to_signed(-23, 8),
    to_signed(-19, 8),
    to_signed(-15, 8),
    to_signed(-10, 8),
    to_signed(-3, 8),
    to_signed(4, 8),
    to_signed(8, 8),
    to_signed(5, 8),
    to_signed(-3, 8),
    to_signed(-12, 8),
    to_signed(-18, 8),
    to_signed(-22, 8),
    to_signed(-22, 8),
    to_signed(-20, 8),
    to_signed(-15, 8),
    to_signed(-8, 8),
    to_signed(2, 8),
    to_signed(12, 8),
    to_signed(21, 8),
    to_signed(28, 8),
    to_signed(34, 8),
    to_signed(40, 8),
    to_signed(43, 8),
    to_signed(40, 8),
    to_signed(34, 8),
    to_signed(27, 8),
    to_signed(20, 8),
    to_signed(14, 8),
    to_signed(8, 8),
    to_signed(4, 8),
    to_signed(6, 8),
    to_signed(14, 8),
    to_signed(27, 8),
    to_signed(41, 8),
    to_signed(52, 8),
    to_signed(59, 8),
    to_signed(62, 8),
    to_signed(60, 8),
    to_signed(51, 8),
    to_signed(35, 8),
    to_signed(15, 8),
    to_signed(-9, 8),
    to_signed(-36, 8),
    to_signed(-64, 8),
    to_signed(-84, 8),
    to_signed(-89, 8),
    to_signed(-77, 8),
    to_signed(-51, 8),
    to_signed(-22, 8),
    to_signed(1, 8),
    to_signed(15, 8),
    to_signed(18, 8),
    to_signed(10, 8),
    to_signed(-9, 8),
    to_signed(-34, 8),
    to_signed(-56, 8),
    to_signed(-67, 8),
    to_signed(-65, 8),
    to_signed(-55, 8),
    to_signed(-41, 8),
    to_signed(-24, 8),
    to_signed(-3, 8),
    to_signed(18, 8),
    to_signed(35, 8),
    to_signed(42, 8),
    to_signed(38, 8),
    to_signed(28, 8),
    to_signed(16, 8),
    to_signed(4, 8),
    to_signed(-9, 8),
    to_signed(-22, 8),
    to_signed(-33, 8),
    to_signed(-40, 8),
    to_signed(-41, 8),
    to_signed(-36, 8),
    to_signed(-29, 8),
    to_signed(-19, 8),
    to_signed(-9, 8),
    to_signed(0, 8),
    to_signed(4, 8),
    to_signed(2, 8),
    to_signed(-5, 8),
    to_signed(-14, 8),
    to_signed(-22, 8),
    to_signed(-25, 8),
    to_signed(-23, 8),
    to_signed(-18, 8),
    to_signed(-13, 8),
    to_signed(-9, 8),
    to_signed(-2, 8),
    to_signed(7, 8),
    to_signed(16, 8),
    to_signed(25, 8),
    to_signed(34, 8),
    to_signed(43, 8),
    to_signed(48, 8),
    to_signed(49, 8),
    to_signed(45, 8),
    to_signed(38, 8),
    to_signed(30, 8),
    to_signed(24, 8),
    to_signed(19, 8),
    to_signed(15, 8),
    to_signed(15, 8),
    to_signed(20, 8),
    to_signed(31, 8),
    to_signed(45, 8),
    to_signed(57, 8),
    to_signed(66, 8),
    to_signed(71, 8),
    to_signed(70, 8),
    to_signed(62, 8),
    to_signed(45, 8),
    to_signed(22, 8),
    to_signed(-6, 8),
    to_signed(-37, 8),
    to_signed(-67, 8),
    to_signed(-88, 8),
    to_signed(-95, 8),
    to_signed(-85, 8),
    to_signed(-62, 8),
    to_signed(-34, 8),
    to_signed(-11, 8),
    to_signed(2, 8),
    to_signed(6, 8),
    to_signed(1, 8),
    to_signed(-14, 8),
    to_signed(-35, 8),
    to_signed(-55, 8),
    to_signed(-67, 8),
    to_signed(-67, 8),
    to_signed(-58, 8),
    to_signed(-45, 8),
    to_signed(-29, 8),
    to_signed(-10, 8),
    to_signed(10, 8),
    to_signed(27, 8),
    to_signed(36, 8),
    to_signed(35, 8),
    to_signed(28, 8),
    to_signed(19, 8),
    to_signed(9, 8),
    to_signed(-2, 8),
    to_signed(-15, 8),
    to_signed(-29, 8),
    to_signed(-39, 8),
    to_signed(-43, 8),
    to_signed(-41, 8),
    to_signed(-34, 8),
    to_signed(-22, 8),
    to_signed(-10, 8),
    to_signed(2, 8),
    to_signed(11, 8),
    to_signed(14, 8),
    to_signed(9, 8),
    to_signed(1, 8),
    to_signed(-8, 8),
    to_signed(-14, 8),
    to_signed(-15, 8),
    to_signed(-13, 8),
    to_signed(-9, 8),
    to_signed(-5, 8),
    to_signed(0, 8),
    to_signed(8, 8),
    to_signed(18, 8),
    to_signed(29, 8),
    to_signed(39, 8),
    to_signed(47, 8),
    to_signed(52, 8),
    to_signed(53, 8),
    to_signed(48, 8),
    to_signed(41, 8),
    to_signed(33, 8),
    to_signed(25, 8),
    to_signed(18, 8),
    to_signed(15, 8),
    to_signed(15, 8),
    to_signed(19, 8),
    to_signed(28, 8),
    to_signed(39, 8),
    to_signed(50, 8),
    to_signed(57, 8),
    to_signed(60, 8),
    to_signed(61, 8),
    to_signed(56, 8),
    to_signed(43, 8),
    to_signed(23, 8),
    to_signed(-3, 8),
    to_signed(-35, 8),
    to_signed(-69, 8),
    to_signed(-94, 8),
    to_signed(-103, 8),
    to_signed(-94, 8),
    to_signed(-71, 8),
    to_signed(-41, 8),
    to_signed(-13, 8),
    to_signed(6, 8),
    to_signed(12, 8),
    to_signed(6, 8),
    to_signed(-10, 8),
    to_signed(-33, 8),
    to_signed(-55, 8),
    to_signed(-69, 8),
    to_signed(-70, 8),
    to_signed(-62, 8),
    to_signed(-49, 8),
    to_signed(-33, 8),
    to_signed(-14, 8),
    to_signed(6, 8),
    to_signed(21, 8),
    to_signed(31, 8),
    to_signed(32, 8),
    to_signed(28, 8),
    to_signed(20, 8),
    to_signed(12, 8),
    to_signed(2, 8),
    to_signed(-10, 8),
    to_signed(-23, 8),
    to_signed(-32, 8),
    to_signed(-35, 8),
    to_signed(-32, 8),
    to_signed(-24, 8),
    to_signed(-13, 8),
    to_signed(-1, 8),
    to_signed(9, 8),
    to_signed(15, 8),
    to_signed(13, 8),
    to_signed(6, 8),
    to_signed(-3, 8),
    to_signed(-11, 8),
    to_signed(-14, 8),
    to_signed(-12, 8),
    to_signed(-8, 8),
    to_signed(-3, 8),
    to_signed(0, 8),
    to_signed(4, 8),
    to_signed(10, 8),
    to_signed(15, 8),
    to_signed(22, 8),
    to_signed(29, 8),
    to_signed(37, 8),
    to_signed(42, 8),
    to_signed(43, 8),
    to_signed(42, 8),
    to_signed(38, 8),
    to_signed(32, 8),
    to_signed(24, 8),
    to_signed(17, 8),
    to_signed(12, 8),
    to_signed(11, 8),
    to_signed(16, 8),
    to_signed(25, 8),
    to_signed(37, 8),
    to_signed(49, 8),
    to_signed(57, 8),
    to_signed(62, 8),
    to_signed(63, 8),
    to_signed(57, 8),
    to_signed(44, 8),
    to_signed(26, 8),
    to_signed(2, 8),
    to_signed(-28, 8),
    to_signed(-59, 8),
    to_signed(-82, 8),
    to_signed(-91, 8),
    to_signed(-84, 8),
    to_signed(-63, 8),
    to_signed(-36, 8),
    to_signed(-10, 8),
    to_signed(7, 8),
    to_signed(12, 8),
    to_signed(6, 8),
    to_signed(-10, 8),
    to_signed(-33, 8),
    to_signed(-54, 8),
    to_signed(-67, 8),
    to_signed(-68, 8),
    to_signed(-60, 8),
    to_signed(-46, 8),
    to_signed(-28, 8),
    to_signed(-9, 8),
    to_signed(9, 8),
    to_signed(24, 8),
    to_signed(33, 8),
    to_signed(36, 8),
    to_signed(33, 8),
    to_signed(27, 8),
    to_signed(20, 8),
    to_signed(10, 8),
    to_signed(-3, 8),
    to_signed(-17, 8),
    to_signed(-28, 8),
    to_signed(-33, 8),
    to_signed(-33, 8),
    to_signed(-28, 8),
    to_signed(-18, 8),
    to_signed(-6, 8),
    to_signed(5, 8),
    to_signed(11, 8),
    to_signed(10, 8),
    to_signed(2, 8),
    to_signed(-10, 8),
    to_signed(-18, 8),
    to_signed(-21, 8),
    to_signed(-19, 8),
    to_signed(-14, 8),
    to_signed(-9, 8),
    to_signed(-5, 8),
    to_signed(-1, 8),
    to_signed(4, 8),
    to_signed(9, 8),
    to_signed(14, 8),
    to_signed(19, 8),
    to_signed(26, 8),
    to_signed(34, 8),
    to_signed(40, 8),
    to_signed(40, 8),
    to_signed(35, 8),
    to_signed(26, 8),
    to_signed(16, 8),
    to_signed(6, 8),
    to_signed(1, 8),
    to_signed(0, 8),
    to_signed(6, 8),
    to_signed(17, 8),
    to_signed(30, 8),
    to_signed(43, 8),
    to_signed(53, 8),
    to_signed(59, 8),
    to_signed(61, 8),
    to_signed(58, 8),
    to_signed(48, 8),
    to_signed(31, 8),
    to_signed(9, 8),
    to_signed(-19, 8),
    to_signed(-51, 8),
    to_signed(-79, 8),
    to_signed(-95, 8),
    to_signed(-92, 8),
    to_signed(-72, 8),
    to_signed(-42, 8),
    to_signed(-12, 8),
    to_signed(11, 8),
    to_signed(21, 8),
    to_signed(19, 8),
    to_signed(4, 8),
    to_signed(-18, 8),
    to_signed(-42, 8),
    to_signed(-60, 8),
    to_signed(-67, 8),
    to_signed(-62, 8),
    to_signed(-50, 8),
    to_signed(-33, 8),
    to_signed(-12, 8),
    to_signed(9, 8),
    to_signed(26, 8),
    to_signed(35, 8),
    to_signed(37, 8),
    to_signed(34, 8),
    to_signed(28, 8),
    to_signed(19, 8),
    to_signed(8, 8),
    to_signed(-5, 8),
    to_signed(-17, 8),
    to_signed(-26, 8),
    to_signed(-30, 8),
    to_signed(-30, 8),
    to_signed(-26, 8),
    to_signed(-20, 8),
    to_signed(-12, 8),
    to_signed(-3, 8),
    to_signed(1, 8),
    to_signed(1, 8),
    to_signed(-5, 8),
    to_signed(-12, 8),
    to_signed(-17, 8),
    to_signed(-19, 8),
    to_signed(-15, 8),
    to_signed(-9, 8),
    to_signed(-5, 8),
    to_signed(-4, 8),
    to_signed(-4, 8),
    to_signed(-1, 8),
    to_signed(2, 8),
    to_signed(6, 8),
    to_signed(11, 8),
    to_signed(21, 8),
    to_signed(34, 8),
    to_signed(45, 8),
    to_signed(52, 8),
    to_signed(52, 8),
    to_signed(46, 8),
    to_signed(34, 8),
    to_signed(22, 8),
    to_signed(13, 8),
    to_signed(9, 8),
    to_signed(10, 8),
    to_signed(20, 8),
    to_signed(33, 8),
    to_signed(47, 8),
    to_signed(56, 8),
    to_signed(64, 8),
    to_signed(70, 8),
    to_signed(70, 8),
    to_signed(60, 8),
    to_signed(43, 8),
    to_signed(20, 8),
    to_signed(-9, 8),
    to_signed(-42, 8),
    to_signed(-73, 8),
    to_signed(-94, 8),
    to_signed(-97, 8),
    to_signed(-80, 8),
    to_signed(-50, 8),
    to_signed(-17, 8),
    to_signed(8, 8),
    to_signed(22, 8),
    to_signed(23, 8),
    to_signed(13, 8),
    to_signed(-8, 8),
    to_signed(-34, 8),
    to_signed(-56, 8),
    to_signed(-68, 8),
    to_signed(-68, 8),
    to_signed(-60, 8),
    to_signed(-45, 8),
    to_signed(-24, 8),
    to_signed(-2, 8),
    to_signed(18, 8),
    to_signed(31, 8),
    to_signed(37, 8),
    to_signed(35, 8),
    to_signed(29, 8),
    to_signed(20, 8),
    to_signed(8, 8),
    to_signed(-6, 8),
    to_signed(-21, 8),
    to_signed(-33, 8),
    to_signed(-39, 8),
    to_signed(-39, 8),
    to_signed(-33, 8),
    to_signed(-25, 8),
    to_signed(-14, 8),
    to_signed(-4, 8),
    to_signed(3, 8),
    to_signed(5, 8),
    to_signed(1, 8),
    to_signed(-8, 8),
    to_signed(-19, 8),
    to_signed(-25, 8),
    to_signed(-25, 8),
    to_signed(-19, 8),
    to_signed(-12, 8),
    to_signed(-6, 8),
    to_signed(-1, 8),
    to_signed(4, 8),
    to_signed(10, 8),
    to_signed(17, 8),
    to_signed(23, 8),
    to_signed(31, 8),
    to_signed(41, 8),
    to_signed(50, 8),
    to_signed(55, 8),
    to_signed(52, 8),
    to_signed(44, 8),
    to_signed(33, 8),
    to_signed(21, 8),
    to_signed(11, 8),
    to_signed(5, 8),
    to_signed(6, 8),
    to_signed(14, 8),
    to_signed(27, 8),
    to_signed(41, 8),
    to_signed(52, 8),
    to_signed(60, 8),
    to_signed(64, 8),
    to_signed(63, 8),
    to_signed(54, 8),
    to_signed(37, 8),
    to_signed(12, 8),
    to_signed(-17, 8),
    to_signed(-50, 8),
    to_signed(-80, 8),
    to_signed(-101, 8),
    to_signed(-103, 8),
    to_signed(-86, 8),
    to_signed(-56, 8),
    to_signed(-24, 8),
    to_signed(1, 8),
    to_signed(14, 8),
    to_signed(15, 8),
    to_signed(5, 8),
    to_signed(-15, 8),
    to_signed(-41, 8),
    to_signed(-62, 8),
    to_signed(-73, 8),
    to_signed(-71, 8),
    to_signed(-60, 8),
    to_signed(-43, 8),
    to_signed(-24, 8),
    to_signed(-3, 8),
    to_signed(17, 8),
    to_signed(31, 8),
    to_signed(38, 8),
    to_signed(36, 8),
    to_signed(29, 8),
    to_signed(19, 8),
    to_signed(8, 8),
    to_signed(-4, 8),
    to_signed(-16, 8),
    to_signed(-26, 8),
    to_signed(-33, 8),
    to_signed(-34, 8),
    to_signed(-30, 8),
    to_signed(-22, 8),
    to_signed(-13, 8),
    to_signed(-2, 8),
    to_signed(6, 8),
    to_signed(11, 8),
    to_signed(9, 8),
    to_signed(1, 8),
    to_signed(-9, 8),
    to_signed(-16, 8),
    to_signed(-18, 8),
    to_signed(-14, 8),
    to_signed(-8, 8),
    to_signed(-3, 8),
    to_signed(1, 8),
    to_signed(6, 8),
    to_signed(12, 8),
    to_signed(18, 8),
    to_signed(23, 8),
    to_signed(29, 8),
    to_signed(37, 8),
    to_signed(44, 8),
    to_signed(46, 8),
    to_signed(43, 8),
    to_signed(35, 8),
    to_signed(24, 8),
    to_signed(12, 8),
    to_signed(4, 8),
    to_signed(0, 8),
    to_signed(0, 8),
    to_signed(7, 8),
    to_signed(19, 8),
    to_signed(32, 8),
    to_signed(44, 8),
    to_signed(53, 8),
    to_signed(57, 8),
    to_signed(56, 8),
    to_signed(49, 8),
    to_signed(35, 8),
    to_signed(15, 8),
    to_signed(-10, 8),
    to_signed(-42, 8),
    to_signed(-74, 8),
    to_signed(-98, 8),
    to_signed(-104, 8),
    to_signed(-93, 8),
    to_signed(-68, 8),
    to_signed(-37, 8),
    to_signed(-9, 8),
    to_signed(10, 8),
    to_signed(18, 8),
    to_signed(14, 8),
    to_signed(-3, 8),
    to_signed(-28, 8),
    to_signed(-52, 8),
    to_signed(-65, 8),
    to_signed(-65, 8),
    to_signed(-56, 8),
    to_signed(-40, 8),
    to_signed(-20, 8),
    to_signed(1, 8),
    to_signed(22, 8),
    to_signed(39, 8),
    to_signed(48, 8),
    to_signed(49, 8),
    to_signed(41, 8),
    to_signed(29, 8),
    to_signed(16, 8),
    to_signed(2, 8),
    to_signed(-12, 8),
    to_signed(-23, 8),
    to_signed(-30, 8),
    to_signed(-31, 8),
    to_signed(-27, 8),
    to_signed(-19, 8),
    to_signed(-8, 8),
    to_signed(4, 8),
    to_signed(14, 8),
    to_signed(19, 8),
    to_signed(17, 8),
    to_signed(8, 8),
    to_signed(-3, 8),
    to_signed(-11, 8),
    to_signed(-13, 8),
    to_signed(-10, 8),
    to_signed(-6, 8),
    to_signed(-2, 8),
    to_signed(2, 8),
    to_signed(7, 8),
    to_signed(11, 8),
    to_signed(14, 8),
    to_signed(16, 8),
    to_signed(20, 8),
    to_signed(28, 8),
    to_signed(37, 8),
    to_signed(42, 8),
    to_signed(42, 8),
    to_signed(36, 8),
    to_signed(26, 8),
    to_signed(15, 8),
    to_signed(4, 8),
    to_signed(-2, 8),
    to_signed(-2, 8),
    to_signed(3, 8),
    to_signed(14, 8),
    to_signed(29, 8),
    to_signed(44, 8),
    to_signed(54, 8),
    to_signed(60, 8),
    to_signed(59, 8),
    to_signed(53, 8),
    to_signed(41, 8),
    to_signed(24, 8),
    to_signed(4, 8),
    to_signed(-23, 8),
    to_signed(-52, 8),
    to_signed(-77, 8),
    to_signed(-89, 8),
    to_signed(-83, 8),
    to_signed(-62, 8),
    to_signed(-35, 8),
    to_signed(-7, 8),
    to_signed(12, 8),
    to_signed(21, 8),
    to_signed(20, 8),
    to_signed(7, 8),
    to_signed(-15, 8),
    to_signed(-38, 8),
    to_signed(-52, 8),
    to_signed(-54, 8),
    to_signed(-47, 8),
    to_signed(-33, 8),
    to_signed(-17, 8),
    to_signed(1, 8),
    to_signed(20, 8),
    to_signed(37, 8),
    to_signed(47, 8),
    to_signed(49, 8),
    to_signed(43, 8),
    to_signed(34, 8),
    to_signed(24, 8),
    to_signed(13, 8),
    to_signed(0, 8),
    to_signed(-12, 8),
    to_signed(-21, 8),
    to_signed(-23, 8),
    to_signed(-22, 8),
    to_signed(-18, 8),
    to_signed(-12, 8),
    to_signed(-5, 8),
    to_signed(3, 8),
    to_signed(9, 8),
    to_signed(8, 8),
    to_signed(2, 8),
    to_signed(-7, 8),
    to_signed(-12, 8),
    to_signed(-14, 8),
    to_signed(-13, 8),
    to_signed(-11, 8),
    to_signed(-9, 8),
    to_signed(-7, 8),
    to_signed(-5, 8),
    to_signed(-1, 8),
    to_signed(2, 8),
    to_signed(6, 8),
    to_signed(12, 8),
    to_signed(21, 8),
    to_signed(33, 8),
    to_signed(42, 8),
    to_signed(46, 8),
    to_signed(42, 8),
    to_signed(32, 8),
    to_signed(20, 8),
    to_signed(9, 8),
    to_signed(2, 8),
    to_signed(-1, 8),
    to_signed(3, 8),
    to_signed(15, 8),
    to_signed(33, 8),
    to_signed(51, 8),
    to_signed(63, 8),
    to_signed(67, 8),
    to_signed(66, 8),
    to_signed(60, 8),
    to_signed(49, 8),
    to_signed(34, 8),
    to_signed(14, 8),
    to_signed(-11, 8),
    to_signed(-40, 8),
    to_signed(-67, 8),
    to_signed(-82, 8),
    to_signed(-83, 8),
    to_signed(-68, 8),
    to_signed(-42, 8),
    to_signed(-14, 8),
    to_signed(6, 8),
    to_signed(16, 8),
    to_signed(16, 8),
    to_signed(6, 8),
    to_signed(-14, 8),
    to_signed(-39, 8),
    to_signed(-57, 8),
    to_signed(-63, 8),
    to_signed(-57, 8),
    to_signed(-42, 8),
    to_signed(-23, 8),
    to_signed(0, 8),
    to_signed(23, 8),
    to_signed(43, 8),
    to_signed(54, 8),
    to_signed(54, 8),
    to_signed(46, 8),
    to_signed(35, 8),
    to_signed(24, 8),
    to_signed(12, 8),
    to_signed(-3, 8),
    to_signed(-16, 8),
    to_signed(-25, 8),
    to_signed(-28, 8),
    to_signed(-29, 8),
    to_signed(-27, 8),
    to_signed(-23, 8),
    to_signed(-17, 8),
    to_signed(-11, 8),
    to_signed(-5, 8),
    to_signed(-2, 8),
    to_signed(-2, 8),
    to_signed(-5, 8),
    to_signed(-8, 8),
    to_signed(-10, 8),
    to_signed(-12, 8),
    to_signed(-12, 8),
    to_signed(-10, 8),
    to_signed(-7, 8),
    to_signed(-5, 8),
    to_signed(-1, 8),
    to_signed(6, 8),
    to_signed(15, 8),
    to_signed(22, 8),
    to_signed(29, 8),
    to_signed(37, 8),
    to_signed(44, 8),
    to_signed(46, 8),
    to_signed(42, 8),
    to_signed(33, 8),
    to_signed(23, 8),
    to_signed(14, 8),
    to_signed(7, 8),
    to_signed(4, 8),
    to_signed(5, 8),
    to_signed(13, 8),
    to_signed(28, 8),
    to_signed(44, 8),
    to_signed(55, 8),
    to_signed(58, 8),
    to_signed(56, 8),
    to_signed(52, 8),
    to_signed(45, 8),
    to_signed(32, 8),
    to_signed(12, 8),
    to_signed(-14, 8),
    to_signed(-44, 8),
    to_signed(-73, 8),
    to_signed(-92, 8),
    to_signed(-94, 8),
    to_signed(-79, 8),
    to_signed(-55, 8),
    to_signed(-29, 8),
    to_signed(-8, 8),
    to_signed(5, 8),
    to_signed(8, 8),
    to_signed(1, 8),
    to_signed(-15, 8),
    to_signed(-36, 8),
    to_signed(-52, 8),
    to_signed(-57, 8),
    to_signed(-51, 8),
    to_signed(-40, 8),
    to_signed(-26, 8),
    to_signed(-7, 8),
    to_signed(15, 8),
    to_signed(34, 8),
    to_signed(45, 8),
    to_signed(46, 8),
    to_signed(42, 8),
    to_signed(35, 8),
    to_signed(26, 8),
    to_signed(14, 8),
    to_signed(0, 8),
    to_signed(-13, 8),
    to_signed(-24, 8),
    to_signed(-29, 8),
    to_signed(-32, 8),
    to_signed(-32, 8),
    to_signed(-30, 8),
    to_signed(-23, 8),
    to_signed(-15, 8),
    to_signed(-9, 8),
    to_signed(-6, 8),
    to_signed(-4, 8),
    to_signed(-3, 8),
    to_signed(-4, 8),
    to_signed(-7, 8),
    to_signed(-11, 8),
    to_signed(-13, 8),
    to_signed(-13, 8),
    to_signed(-13, 8),
    to_signed(-12, 8),
    to_signed(-8, 8),
    to_signed(-3, 8),
    to_signed(5, 8),
    to_signed(14, 8),
    to_signed(24, 8),
    to_signed(34, 8),
    to_signed(42, 8),
    to_signed(46, 8),
    to_signed(43, 8),
    to_signed(35, 8),
    to_signed(24, 8),
    to_signed(13, 8),
    to_signed(3, 8),
    to_signed(-3, 8),
    to_signed(-3, 8),
    to_signed(6, 8),
    to_signed(22, 8),
    to_signed(40, 8),
    to_signed(51, 8),
    to_signed(56, 8),
    to_signed(55, 8),
    to_signed(50, 8),
    to_signed(38, 8),
    to_signed(19, 8),
    to_signed(-4, 8),
    to_signed(-31, 8),
    to_signed(-59, 8),
    to_signed(-83, 8),
    to_signed(-95, 8),
    to_signed(-89, 8),
    to_signed(-69, 8),
    to_signed(-42, 8),
    to_signed(-16, 8),
    to_signed(1, 8),
    to_signed(8, 8),
    to_signed(7, 8),
    to_signed(-2, 8),
    to_signed(-19, 8),
    to_signed(-38, 8),
    to_signed(-51, 8),
    to_signed(-51, 8),
    to_signed(-42, 8),
    to_signed(-30, 8),
    to_signed(-17, 8),
    to_signed(1, 8),
    to_signed(20, 8),
    to_signed(36, 8),
    to_signed(45, 8),
    to_signed(46, 8),
    to_signed(41, 8),
    to_signed(31, 8),
    to_signed(20, 8),
    to_signed(8, 8),
    to_signed(-5, 8),
    to_signed(-16, 8),
    to_signed(-24, 8),
    to_signed(-28, 8),
    to_signed(-28, 8),
    to_signed(-26, 8),
    to_signed(-21, 8),
    to_signed(-14, 8),
    to_signed(-9, 8),
    to_signed(-8, 8),
    to_signed(-10, 8),
    to_signed(-11, 8),
    to_signed(-12, 8),
    to_signed(-15, 8),
    to_signed(-16, 8),
    to_signed(-15, 8),
    to_signed(-13, 8),
    to_signed(-11, 8),
    to_signed(-11, 8),
    to_signed(-10, 8),
    to_signed(-7, 8),
    to_signed(-1, 8),
    to_signed(6, 8),
    to_signed(15, 8),
    to_signed(25, 8),
    to_signed(36, 8),
    to_signed(45, 8),
    to_signed(48, 8),
    to_signed(42, 8),
    to_signed(31, 8),
    to_signed(19, 8),
    to_signed(9, 8),
    to_signed(1, 8),
    to_signed(-4, 8),
    to_signed(-2, 8),
    to_signed(11, 8),
    to_signed(28, 8),
    to_signed(45, 8),
    to_signed(56, 8),
    to_signed(60, 8),
    to_signed(59, 8),
    to_signed(51, 8),
    to_signed(38, 8),
    to_signed(18, 8),
    to_signed(-6, 8),
    to_signed(-33, 8),
    to_signed(-60, 8),
    to_signed(-80, 8),
    to_signed(-88, 8),
    to_signed(-79, 8),
    to_signed(-56, 8),
    to_signed(-27, 8),
    to_signed(-3, 8),
    to_signed(13, 8),
    to_signed(18, 8),
    to_signed(13, 8),
    to_signed(-2, 8),
    to_signed(-24, 8),
    to_signed(-46, 8),
    to_signed(-57, 8),
    to_signed(-55, 8),
    to_signed(-43, 8),
    to_signed(-28, 8),
    to_signed(-10, 8),
    to_signed(11, 8),
    to_signed(31, 8),
    to_signed(45, 8),
    to_signed(49, 8),
    to_signed(45, 8),
    to_signed(36, 8),
    to_signed(24, 8),
    to_signed(11, 8),
    to_signed(-2, 8),
    to_signed(-12, 8),
    to_signed(-19, 8),
    to_signed(-23, 8),
    to_signed(-26, 8),
    to_signed(-28, 8),
    to_signed(-27, 8),
    to_signed(-21, 8),
    to_signed(-14, 8),
    to_signed(-10, 8),
    to_signed(-9, 8),
    to_signed(-11, 8),
    to_signed(-11, 8),
    to_signed(-13, 8),
    to_signed(-16, 8),
    to_signed(-17, 8),
    to_signed(-14, 8),
    to_signed(-10, 8),
    to_signed(-6, 8),
    to_signed(-4, 8),
    to_signed(-3, 8),
    to_signed(1, 8),
    to_signed(7, 8),
    to_signed(15, 8),
    to_signed(23, 8),
    to_signed(32, 8),
    to_signed(40, 8),
    to_signed(46, 8),
    to_signed(45, 8),
    to_signed(37, 8),
    to_signed(26, 8),
    to_signed(14, 8),
    to_signed(6, 8),
    to_signed(0, 8),
    to_signed(-2, 8),
    to_signed(3, 8),
    to_signed(17, 8),
    to_signed(36, 8),
    to_signed(51, 8),
    to_signed(61, 8),
    to_signed(63, 8),
    to_signed(60, 8),
    to_signed(52, 8),
    to_signed(37, 8),
    to_signed(18, 8),
    to_signed(-4, 8),
    to_signed(-28, 8),
    to_signed(-53, 8),
    to_signed(-73, 8),
    to_signed(-82, 8),
    to_signed(-76, 8),
    to_signed(-57, 8),
    to_signed(-33, 8),
    to_signed(-11, 8),
    to_signed(4, 8),
    to_signed(13, 8),
    to_signed(12, 8),
    to_signed(-1, 8),
    to_signed(-23, 8),
    to_signed(-45, 8),
    to_signed(-58, 8),
    to_signed(-59, 8),
    to_signed(-52, 8),
    to_signed(-41, 8),
    to_signed(-25, 8),
    to_signed(-3, 8),
    to_signed(20, 8),
    to_signed(38, 8),
    to_signed(46, 8),
    to_signed(45, 8),
    to_signed(37, 8),
    to_signed(25, 8),
    to_signed(10, 8),
    to_signed(-7, 8),
    to_signed(-20, 8),
    to_signed(-29, 8),
    to_signed(-33, 8),
    to_signed(-35, 8),
    to_signed(-35, 8),
    to_signed(-32, 8),
    to_signed(-24, 8),
    to_signed(-15, 8),
    to_signed(-8, 8),
    to_signed(-4, 8),
    to_signed(-4, 8),
    to_signed(-5, 8),
    to_signed(-8, 8),
    to_signed(-12, 8),
    to_signed(-14, 8),
    to_signed(-11, 8),
    to_signed(-6, 8),
    to_signed(0, 8),
    to_signed(2, 8),
    to_signed(3, 8),
    to_signed(5, 8),
    to_signed(8, 8),
    to_signed(13, 8),
    to_signed(20, 8),
    to_signed(29, 8),
    to_signed(39, 8),
    to_signed(47, 8),
    to_signed(49, 8),
    to_signed(43, 8),
    to_signed(33, 8),
    to_signed(21, 8),
    to_signed(10, 8),
    to_signed(1, 8),
    to_signed(-3, 8),
    to_signed(-1, 8),
    to_signed(10, 8),
    to_signed(27, 8),
    to_signed(45, 8),
    to_signed(56, 8),
    to_signed(61, 8),
    to_signed(60, 8),
    to_signed(53, 8),
    to_signed(39, 8),
    to_signed(19, 8),
    to_signed(-4, 8),
    to_signed(-31, 8),
    to_signed(-58, 8),
    to_signed(-79, 8),
    to_signed(-87, 8),
    to_signed(-78, 8),
    to_signed(-58, 8),
    to_signed(-34, 8),
    to_signed(-13, 8),
    to_signed(4, 8),
    to_signed(13, 8),
    to_signed(13, 8),
    to_signed(1, 8),
    to_signed(-19, 8),
    to_signed(-41, 8),
    to_signed(-55, 8),
    to_signed(-58, 8),
    to_signed(-54, 8),
    to_signed(-46, 8),
    to_signed(-31, 8),
    to_signed(-8, 8),
    to_signed(17, 8),
    to_signed(37, 8),
    to_signed(48, 8),
    to_signed(51, 8),
    to_signed(47, 8),
    to_signed(36, 8),
    to_signed(21, 8),
    to_signed(6, 8),
    to_signed(-8, 8),
    to_signed(-19, 8),
    to_signed(-25, 8),
    to_signed(-26, 8),
    to_signed(-26, 8),
    to_signed(-25, 8),
    to_signed(-20, 8),
    to_signed(-12, 8),
    to_signed(-4, 8),
    to_signed(0, 8),
    to_signed(2, 8),
    to_signed(1, 8),
    to_signed(-2, 8),
    to_signed(-9, 8),
    to_signed(-15, 8),
    to_signed(-16, 8),
    to_signed(-15, 8),
    to_signed(-12, 8),
    to_signed(-9, 8),
    to_signed(-4, 8),
    to_signed(3, 8),
    to_signed(8, 8),
    to_signed(16, 8),
    to_signed(25, 8),
    to_signed(35, 8),
    to_signed(43, 8),
    to_signed(49, 8),
    to_signed(51, 8),
    to_signed(46, 8),
    to_signed(36, 8),
    to_signed(26, 8),
    to_signed(18, 8),
    to_signed(12, 8),
    to_signed(9, 8),
    to_signed(12, 8),
    to_signed(21, 8),
    to_signed(34, 8),
    to_signed(45, 8),
    to_signed(54, 8),
    to_signed(60, 8),
    to_signed(60, 8),
    to_signed(53, 8),
    to_signed(38, 8),
    to_signed(17, 8),
    to_signed(-9, 8),
    to_signed(-40, 8),
    to_signed(-69, 8),
    to_signed(-87, 8),
    to_signed(-89, 8),
    to_signed(-74, 8),
    to_signed(-50, 8),
    to_signed(-25, 8),
    to_signed(-5, 8),
    to_signed(7, 8),
    to_signed(10, 8),
    to_signed(5, 8),
    to_signed(-9, 8),
    to_signed(-28, 8),
    to_signed(-45, 8),
    to_signed(-53, 8),
    to_signed(-51, 8),
    to_signed(-43, 8),
    to_signed(-32, 8),
    to_signed(-15, 8),
    to_signed(7, 8),
    to_signed(28, 8),
    to_signed(42, 8),
    to_signed(49, 8),
    to_signed(49, 8),
    to_signed(42, 8),
    to_signed(31, 8),
    to_signed(19, 8),
    to_signed(6, 8),
    to_signed(-6, 8),
    to_signed(-18, 8),
    to_signed(-23, 8),
    to_signed(-24, 8),
    to_signed(-24, 8),
    to_signed(-24, 8),
    to_signed(-22, 8),
    to_signed(-17, 8),
    to_signed(-11, 8),
    to_signed(-6, 8),
    to_signed(-2, 8),
    to_signed(0, 8),
    to_signed(-3, 8),
    to_signed(-8, 8),
    to_signed(-10, 8),
    to_signed(-8, 8),
    to_signed(-6, 8),
    to_signed(-6, 8),
    to_signed(-5, 8),
    to_signed(-1, 8),
    to_signed(4, 8),
    to_signed(8, 8),
    to_signed(15, 8),
    to_signed(25, 8),
    to_signed(34, 8),
    to_signed(40, 8),
    to_signed(44, 8),
    to_signed(44, 8),
    to_signed(36, 8),
    to_signed(23, 8),
    to_signed(13, 8),
    to_signed(7, 8),
    to_signed(3, 8),
    to_signed(4, 8),
    to_signed(13, 8),
    to_signed(28, 8),
    to_signed(43, 8),
    to_signed(53, 8),
    to_signed(61, 8),
    to_signed(63, 8),
    to_signed(58, 8),
    to_signed(43, 8),
    to_signed(21, 8),
    to_signed(-5, 8),
    to_signed(-35, 8),
    to_signed(-66, 8),
    to_signed(-88, 8),
    to_signed(-93, 8),
    to_signed(-83, 8),
    to_signed(-62, 8),
    to_signed(-36, 8),
    to_signed(-15, 8),
    to_signed(-4, 8),
    to_signed(-4, 8),
    to_signed(-10, 8),
    to_signed(-22, 8),
    to_signed(-36, 8),
    to_signed(-49, 8),
    to_signed(-52, 8),
    to_signed(-45, 8),
    to_signed(-34, 8),
    to_signed(-23, 8),
    to_signed(-9, 8),
    to_signed(7, 8),
    to_signed(23, 8),
    to_signed(34, 8),
    to_signed(41, 8),
    to_signed(44, 8),
    to_signed(42, 8),
    to_signed(34, 8),
    to_signed(23, 8),
    to_signed(13, 8),
    to_signed(2, 8),
    to_signed(-10, 8),
    to_signed(-22, 8),
    to_signed(-29, 8),
    to_signed(-30, 8),
    to_signed(-27, 8),
    to_signed(-21, 8),
    to_signed(-14, 8),
    to_signed(-11, 8),
    to_signed(-10, 8),
    to_signed(-9, 8),
    to_signed(-7, 8),
    to_signed(-8, 8),
    to_signed(-11, 8),
    to_signed(-13, 8),
    to_signed(-10, 8),
    to_signed(-4, 8),
    to_signed(1, 8),
    to_signed(2, 8),
    to_signed(2, 8),
    to_signed(1, 8),
    to_signed(1, 8),
    to_signed(3, 8),
    to_signed(9, 8),
    to_signed(18, 8),
    to_signed(27, 8),
    to_signed(34, 8),
    to_signed(38, 8),
    to_signed(37, 8),
    to_signed(28, 8),
    to_signed(15, 8),
    to_signed(5, 8),
    to_signed(-1, 8),
    to_signed(-1, 8),
    to_signed(7, 8),
    to_signed(22, 8),
    to_signed(39, 8),
    to_signed(54, 8),
    to_signed(62, 8),
    to_signed(66, 8),
    to_signed(63, 8),
    to_signed(50, 8),
    to_signed(30, 8),
    to_signed(5, 8),
    to_signed(-22, 8),
    to_signed(-51, 8),
    to_signed(-79, 8),
    to_signed(-95, 8),
    to_signed(-92, 8),
    to_signed(-71, 8),
    to_signed(-43, 8),
    to_signed(-18, 8),
    to_signed(-2, 8),
    to_signed(3, 8),
    to_signed(-1, 8),
    to_signed(-10, 8),
    to_signed(-24, 8),
    to_signed(-41, 8),
    to_signed(-52, 8),
    to_signed(-49, 8),
    to_signed(-37, 8),
    to_signed(-23, 8),
    to_signed(-10, 8),
    to_signed(5, 8),
    to_signed(21, 8),
    to_signed(33, 8),
    to_signed(37, 8),
    to_signed(34, 8),
    to_signed(29, 8),
    to_signed(22, 8),
    to_signed(15, 8),
    to_signed(8, 8),
    to_signed(1, 8),
    to_signed(-7, 8),
    to_signed(-15, 8),
    to_signed(-23, 8),
    to_signed(-29, 8),
    to_signed(-33, 8),
    to_signed(-32, 8),
    to_signed(-24, 8),
    to_signed(-15, 8),
    to_signed(-11, 8),
    to_signed(-11, 8),
    to_signed(-11, 8),
    to_signed(-11, 8),
    to_signed(-12, 8),
    to_signed(-14, 8),
    to_signed(-13, 8),
    to_signed(-9, 8),
    to_signed(-3, 8),
    to_signed(1, 8),
    to_signed(3, 8),
    to_signed(2, 8),
    to_signed(0, 8),
    to_signed(-1, 8),
    to_signed(1, 8),
    to_signed(8, 8),
    to_signed(17, 8),
    to_signed(27, 8),
    to_signed(35, 8),
    to_signed(38, 8),
    to_signed(35, 8),
    to_signed(28, 8),
    to_signed(19, 8),
    to_signed(10, 8),
    to_signed(2, 8),
    to_signed(1, 8),
    to_signed(9, 8),
    to_signed(25, 8),
    to_signed(43, 8),
    to_signed(56, 8),
    to_signed(64, 8),
    to_signed(66, 8),
    to_signed(61, 8),
    to_signed(48, 8),
    to_signed(28, 8),
    to_signed(4, 8),
    to_signed(-22, 8),
    to_signed(-49, 8),
    to_signed(-73, 8),
    to_signed(-89, 8),
    to_signed(-87, 8),
    to_signed(-67, 8),
    to_signed(-37, 8),
    to_signed(-12, 8),
    to_signed(1, 8),
    to_signed(4, 8),
    to_signed(2, 8),
    to_signed(-5, 8),
    to_signed(-17, 8),
    to_signed(-32, 8),
    to_signed(-43, 8),
    to_signed(-46, 8),
    to_signed(-41, 8),
    to_signed(-33, 8),
    to_signed(-24, 8),
    to_signed(-12, 8),
    to_signed(4, 8),
    to_signed(20, 8),
    to_signed(29, 8),
    to_signed(31, 8),
    to_signed(28, 8),
    to_signed(24, 8),
    to_signed(18, 8),
    to_signed(12, 8),
    to_signed(4, 8),
    to_signed(-4, 8),
    to_signed(-14, 8),
    to_signed(-24, 8),
    to_signed(-32, 8),
    to_signed(-34, 8),
    to_signed(-31, 8),
    to_signed(-21, 8),
    to_signed(-9, 8),
    to_signed(0, 8),
    to_signed(2, 8),
    to_signed(-1, 8),
    to_signed(-5, 8),
    to_signed(-9, 8),
    to_signed(-12, 8),
    to_signed(-13, 8),
    to_signed(-9, 8),
    to_signed(-2, 8),
    to_signed(3, 8),
    to_signed(6, 8),
    to_signed(6, 8),
    to_signed(6, 8),
    to_signed(7, 8),
    to_signed(10, 8),
    to_signed(17, 8),
    to_signed(27, 8),
    to_signed(35, 8),
    to_signed(41, 8),
    to_signed(44, 8),
    to_signed(43, 8),
    to_signed(37, 8),
    to_signed(29, 8),
    to_signed(20, 8),
    to_signed(11, 8),
    to_signed(6, 8),
    to_signed(10, 8),
    to_signed(24, 8),
    to_signed(42, 8),
    to_signed(57, 8),
    to_signed(66, 8),
    to_signed(70, 8),
    to_signed(67, 8),
    to_signed(53, 8),
    to_signed(32, 8),
    to_signed(8, 8),
    to_signed(-19, 8),
    to_signed(-47, 8),
    to_signed(-72, 8),
    to_signed(-85, 8),
    to_signed(-81, 8),
    to_signed(-61, 8),
    to_signed(-34, 8),
    to_signed(-10, 8),
    to_signed(4, 8),
    to_signed(7, 8),
    to_signed(3, 8),
    to_signed(-5, 8),
    to_signed(-16, 8),
    to_signed(-29, 8),
    to_signed(-39, 8),
    to_signed(-41, 8),
    to_signed(-39, 8),
    to_signed(-34, 8),
    to_signed(-26, 8),
    to_signed(-15, 8),
    to_signed(0, 8),
    to_signed(15, 8),
    to_signed(26, 8),
    to_signed(32, 8),
    to_signed(34, 8),
    to_signed(32, 8),
    to_signed(27, 8),
    to_signed(19, 8),
    to_signed(9, 8),
    to_signed(-4, 8),
    to_signed(-16, 8),
    to_signed(-27, 8),
    to_signed(-34, 8),
    to_signed(-35, 8),
    to_signed(-29, 8),
    to_signed(-18, 8),
    to_signed(-3, 8),
    to_signed(9, 8),
    to_signed(13, 8),
    to_signed(11, 8),
    to_signed(4, 8),
    to_signed(-3, 8),
    to_signed(-9, 8),
    to_signed(-9, 8),
    to_signed(-4, 8),
    to_signed(4, 8),
    to_signed(9, 8),
    to_signed(11, 8),
    to_signed(12, 8),
    to_signed(11, 8),
    to_signed(11, 8),
    to_signed(14, 8),
    to_signed(21, 8),
    to_signed(30, 8),
    to_signed(38, 8),
    to_signed(42, 8),
    to_signed(43, 8),
    to_signed(41, 8),
    to_signed(35, 8),
    to_signed(27, 8),
    to_signed(18, 8),
    to_signed(10, 8),
    to_signed(6, 8),
    to_signed(10, 8),
    to_signed(22, 8),
    to_signed(38, 8),
    to_signed(51, 8),
    to_signed(61, 8),
    to_signed(66, 8),
    to_signed(61, 8),
    to_signed(46, 8),
    to_signed(23, 8),
    to_signed(-4, 8),
    to_signed(-33, 8),
    to_signed(-62, 8),
    to_signed(-85, 8),
    to_signed(-95, 8),
    to_signed(-86, 8),
    to_signed(-63, 8),
    to_signed(-35, 8),
    to_signed(-10, 8),
    to_signed(6, 8),
    to_signed(11, 8),
    to_signed(6, 8),
    to_signed(-6, 8),
    to_signed(-23, 8),
    to_signed(-39, 8),
    to_signed(-50, 8),
    to_signed(-51, 8),
    to_signed(-47, 8),
    to_signed(-38, 8),
    to_signed(-25, 8),
    to_signed(-7, 8),
    to_signed(10, 8),
    to_signed(22, 8),
    to_signed(28, 8),
    to_signed(29, 8),
    to_signed(26, 8),
    to_signed(21, 8),
    to_signed(13, 8),
    to_signed(3, 8),
    to_signed(-6, 8),
    to_signed(-14, 8),
    to_signed(-21, 8),
    to_signed(-26, 8),
    to_signed(-29, 8),
    to_signed(-27, 8),
    to_signed(-22, 8),
    to_signed(-14, 8),
    to_signed(-4, 8),
    to_signed(3, 8),
    to_signed(7, 8),
    to_signed(7, 8),
    to_signed(2, 8),
    to_signed(-4, 8),
    to_signed(-11, 8),
    to_signed(-11, 8),
    to_signed(-5, 8),
    to_signed(2, 8),
    to_signed(8, 8),
    to_signed(10, 8),
    to_signed(12, 8),
    to_signed(13, 8),
    to_signed(16, 8),
    to_signed(19, 8),
    to_signed(25, 8),
    to_signed(32, 8),
    to_signed(39, 8),
    to_signed(41, 8),
    to_signed(39, 8),
    to_signed(35, 8),
    to_signed(28, 8),
    to_signed(21, 8),
    to_signed(14, 8),
    to_signed(10, 8),
    to_signed(9, 8),
    to_signed(14, 8),
    to_signed(25, 8),
    to_signed(36, 8),
    to_signed(43, 8),
    to_signed(47, 8),
    to_signed(47, 8),
    to_signed(41, 8),
    to_signed(26, 8),
    to_signed(4, 8),
    to_signed(-23, 8),
    to_signed(-51, 8),
    to_signed(-78, 8),
    to_signed(-97, 8),
    to_signed(-101, 8),
    to_signed(-87, 8),
    to_signed(-62, 8),
    to_signed(-36, 8),
    to_signed(-15, 8),
    to_signed(-3, 8),
    to_signed(-1, 8),
    to_signed(-8, 8),
    to_signed(-22, 8),
    to_signed(-38, 8),
    to_signed(-53, 8),
    to_signed(-59, 8),
    to_signed(-55, 8),
    to_signed(-46, 8),
    to_signed(-35, 8),
    to_signed(-20, 8),
    to_signed(1, 8),
    to_signed(19, 8),
    to_signed(29, 8),
    to_signed(31, 8),
    to_signed(29, 8),
    to_signed(26, 8),
    to_signed(22, 8),
    to_signed(17, 8),
    to_signed(11, 8),
    to_signed(4, 8),
    to_signed(-1, 8),
    to_signed(-5, 8),
    to_signed(-9, 8),
    to_signed(-12, 8),
    to_signed(-13, 8),
    to_signed(-10, 8),
    to_signed(-3, 8),
    to_signed(4, 8),
    to_signed(7, 8),
    to_signed(8, 8),
    to_signed(9, 8),
    to_signed(7, 8),
    to_signed(1, 8),
    to_signed(-6, 8),
    to_signed(-8, 8),
    to_signed(-3, 8),
    to_signed(5, 8),
    to_signed(13, 8),
    to_signed(18, 8),
    to_signed(18, 8),
    to_signed(18, 8),
    to_signed(20, 8),
    to_signed(23, 8),
    to_signed(26, 8),
    to_signed(29, 8),
    to_signed(31, 8),
    to_signed(31, 8),
    to_signed(29, 8),
    to_signed(23, 8),
    to_signed(15, 8),
    to_signed(5, 8),
    to_signed(-2, 8),
    to_signed(-6, 8),
    to_signed(-5, 8),
    to_signed(5, 8),
    to_signed(18, 8),
    to_signed(30, 8),
    to_signed(38, 8),
    to_signed(43, 8),
    to_signed(45, 8),
    to_signed(40, 8),
    to_signed(29, 8),
    to_signed(12, 8),
    to_signed(-13, 8),
    to_signed(-42, 8),
    to_signed(-72, 8),
    to_signed(-91, 8),
    to_signed(-93, 8),
    to_signed(-76, 8),
    to_signed(-47, 8),
    to_signed(-18, 8),
    to_signed(3, 8),
    to_signed(14, 8),
    to_signed(16, 8),
    to_signed(7, 8),
    to_signed(-11, 8),
    to_signed(-30, 8),
    to_signed(-45, 8),
    to_signed(-50, 8),
    to_signed(-43, 8),
    to_signed(-32, 8),
    to_signed(-17, 8),
    to_signed(1, 8),
    to_signed(22, 8),
    to_signed(40, 8),
    to_signed(49, 8),
    to_signed(49, 8),
    to_signed(43, 8),
    to_signed(35, 8),
    to_signed(28, 8),
    to_signed(21, 8),
    to_signed(13, 8),
    to_signed(5, 8),
    to_signed(-2, 8),
    to_signed(-8, 8),
    to_signed(-14, 8),
    to_signed(-19, 8),
    to_signed(-22, 8),
    to_signed(-20, 8),
    to_signed(-14, 8),
    to_signed(-7, 8),
    to_signed(-4, 8),
    to_signed(-4, 8),
    to_signed(-4, 8),
    to_signed(-4, 8),
    to_signed(-6, 8),
    to_signed(-10, 8),
    to_signed(-11, 8),
    to_signed(-8, 8),
    to_signed(0, 8),
    to_signed(7, 8),
    to_signed(11, 8),
    to_signed(11, 8),
    to_signed(11, 8),
    to_signed(14, 8),
    to_signed(19, 8),
    to_signed(26, 8),
    to_signed(33, 8),
    to_signed(37, 8),
    to_signed(37, 8),
    to_signed(33, 8),
    to_signed(27, 8),
    to_signed(15, 8),
    to_signed(2, 8),
    to_signed(-8, 8),
    to_signed(-12, 8),
    to_signed(-6, 8),
    to_signed(9, 8),
    to_signed(28, 8),
    to_signed(45, 8),
    to_signed(58, 8),
    to_signed(66, 8),
    to_signed(68, 8),
    to_signed(62, 8),
    to_signed(47, 8),
    to_signed(26, 8),
    to_signed(-1, 8),
    to_signed(-35, 8),
    to_signed(-69, 8),
    to_signed(-91, 8),
    to_signed(-94, 8),
    to_signed(-75, 8),
    to_signed(-45, 8),
    to_signed(-15, 8),
    to_signed(7, 8),
    to_signed(20, 8),
    to_signed(22, 8),
    to_signed(12, 8),
    to_signed(-5, 8),
    to_signed(-25, 8),
    to_signed(-42, 8),
    to_signed(-49, 8),
    to_signed(-46, 8),
    to_signed(-38, 8),
    to_signed(-27, 8),
    to_signed(-10, 8),
    to_signed(10, 8),
    to_signed(27, 8),
    to_signed(38, 8),
    to_signed(40, 8),
    to_signed(35, 8),
    to_signed(27, 8),
    to_signed(17, 8),
    to_signed(7, 8),
    to_signed(-4, 8),
    to_signed(-14, 8),
    to_signed(-22, 8),
    to_signed(-28, 8),
    to_signed(-32, 8),
    to_signed(-35, 8),
    to_signed(-35, 8),
    to_signed(-30, 8),
    to_signed(-22, 8),
    to_signed(-15, 8),
    to_signed(-11, 8),
    to_signed(-11, 8),
    to_signed(-11, 8),
    to_signed(-11, 8),
    to_signed(-12, 8),
    to_signed(-13, 8),
    to_signed(-13, 8),
    to_signed(-11, 8),
    to_signed(-7, 8),
    to_signed(-3, 8),
    to_signed(-1, 8),
    to_signed(0, 8),
    to_signed(3, 8),
    to_signed(9, 8),
    to_signed(20, 8),
    to_signed(33, 8),
    to_signed(44, 8),
    to_signed(51, 8),
    to_signed(50, 8),
    to_signed(44, 8),
    to_signed(34, 8),
    to_signed(22, 8),
    to_signed(9, 8),
    to_signed(-2, 8),
    to_signed(-4, 8),
    to_signed(4, 8),
    to_signed(19, 8),
    to_signed(38, 8),
    to_signed(54, 8),
    to_signed(66, 8),
    to_signed(74, 8),
    to_signed(73, 8),
    to_signed(63, 8),
    to_signed(44, 8),
    to_signed(19, 8),
    to_signed(-12, 8),
    to_signed(-47, 8),
    to_signed(-81, 8),
    to_signed(-102, 8),
    to_signed(-103, 8),
    to_signed(-81, 8),
    to_signed(-49, 8),
    to_signed(-18, 8),
    to_signed(5, 8),
    to_signed(16, 8),
    to_signed(15, 8),
    to_signed(3, 8),
    to_signed(-17, 8),
    to_signed(-38, 8),
    to_signed(-53, 8),
    to_signed(-58, 8),
    to_signed(-54, 8),
    to_signed(-45, 8),
    to_signed(-32, 8),
    to_signed(-17, 8),
    to_signed(1, 8),
    to_signed(16, 8),
    to_signed(24, 8),
    to_signed(27, 8),
    to_signed(24, 8),
    to_signed(18, 8),
    to_signed(13, 8),
    to_signed(4, 8),
    to_signed(-7, 8),
    to_signed(-18, 8),
    to_signed(-26, 8),
    to_signed(-32, 8),
    to_signed(-37, 8),
    to_signed(-38, 8),
    to_signed(-34, 8),
    to_signed(-27, 8),
    to_signed(-18, 8),
    to_signed(-11, 8),
    to_signed(-8, 8),
    to_signed(-9, 8),
    to_signed(-10, 8),
    to_signed(-12, 8),
    to_signed(-14, 8),
    to_signed(-12, 8),
    to_signed(-7, 8),
    to_signed(-1, 8),
    to_signed(5, 8),
    to_signed(10, 8),
    to_signed(12, 8),
    to_signed(13, 8),
    to_signed(16, 8),
    to_signed(22, 8),
    to_signed(31, 8),
    to_signed(43, 8),
    to_signed(57, 8),
    to_signed(65, 8),
    to_signed(64, 8),
    to_signed(56, 8),
    to_signed(43, 8),
    to_signed(28, 8),
    to_signed(12, 8),
    to_signed(0, 8),
    to_signed(-3, 8),
    to_signed(5, 8),
    to_signed(21, 8),
    to_signed(38, 8),
    to_signed(53, 8),
    to_signed(64, 8),
    to_signed(69, 8),
    to_signed(67, 8),
    to_signed(56, 8),
    to_signed(38, 8),
    to_signed(12, 8),
    to_signed(-19, 8),
    to_signed(-50, 8),
    to_signed(-78, 8),
    to_signed(-95, 8),
    to_signed(-95, 8),
    to_signed(-75, 8),
    to_signed(-46, 8),
    to_signed(-20, 8),
    to_signed(-1, 8),
    to_signed(7, 8),
    to_signed(5, 8),
    to_signed(-8, 8),
    to_signed(-26, 8),
    to_signed(-45, 8),
    to_signed(-59, 8),
    to_signed(-65, 8),
    to_signed(-62, 8),
    to_signed(-54, 8),
    to_signed(-42, 8),
    to_signed(-27, 8),
    to_signed(-9, 8),
    to_signed(7, 8),
    to_signed(17, 8),
    to_signed(19, 8),
    to_signed(17, 8),
    to_signed(15, 8),
    to_signed(11, 8),
    to_signed(2, 8),
    to_signed(-9, 8),
    to_signed(-20, 8),
    to_signed(-30, 8),
    to_signed(-37, 8),
    to_signed(-41, 8),
    to_signed(-40, 8),
    to_signed(-35, 8),
    to_signed(-26, 8),
    to_signed(-14, 8),
    to_signed(-6, 8),
    to_signed(-3, 8),
    to_signed(-3, 8),
    to_signed(-4, 8),
    to_signed(-6, 8),
    to_signed(-8, 8),
    to_signed(-7, 8),
    to_signed(-2, 8),
    to_signed(5, 8),
    to_signed(11, 8),
    to_signed(15, 8),
    to_signed(17, 8),
    to_signed(18, 8),
    to_signed(21, 8),
    to_signed(25, 8),
    to_signed(32, 8),
    to_signed(41, 8),
    to_signed(51, 8),
    to_signed(57, 8),
    to_signed(58, 8),
    to_signed(54, 8),
    to_signed(43, 8),
    to_signed(30, 8),
    to_signed(16, 8),
    to_signed(6, 8),
    to_signed(3, 8),
    to_signed(11, 8),
    to_signed(26, 8),
    to_signed(44, 8),
    to_signed(58, 8),
    to_signed(69, 8),
    to_signed(73, 8),
    to_signed(67, 8),
    to_signed(53, 8),
    to_signed(32, 8),
    to_signed(6, 8),
    to_signed(-26, 8),
    to_signed(-57, 8),
    to_signed(-82, 8),
    to_signed(-95, 8),
    to_signed(-92, 8),
    to_signed(-73, 8),
    to_signed(-47, 8),
    to_signed(-24, 8),
    to_signed(-9, 8),
    to_signed(-4, 8),
    to_signed(-10, 8),
    to_signed(-23, 8),
    to_signed(-40, 8),
    to_signed(-54, 8),
    to_signed(-62, 8),
    to_signed(-60, 8),
    to_signed(-53, 8),
    to_signed(-43, 8),
    to_signed(-30, 8),
    to_signed(-14, 8),
    to_signed(3, 8),
    to_signed(16, 8),
    to_signed(24, 8),
    to_signed(23, 8),
    to_signed(18, 8),
    to_signed(14, 8),
    to_signed(11, 8),
    to_signed(5, 8),
    to_signed(-2, 8),
    to_signed(-9, 8),
    to_signed(-15, 8),
    to_signed(-21, 8),
    to_signed(-25, 8),
    to_signed(-26, 8),
    to_signed(-24, 8),
    to_signed(-18, 8),
    to_signed(-11, 8),
    to_signed(-5, 8),
    to_signed(-2, 8),
    to_signed(-2, 8),
    to_signed(-1, 8),
    to_signed(-1, 8),
    to_signed(2, 8),
    to_signed(6, 8),
    to_signed(13, 8),
    to_signed(18, 8),
    to_signed(20, 8),
    to_signed(20, 8),
    to_signed(17, 8),
    to_signed(14, 8),
    to_signed(14, 8),
    to_signed(18, 8),
    to_signed(26, 8),
    to_signed(38, 8),
    to_signed(50, 8),
    to_signed(58, 8),
    to_signed(60, 8),
    to_signed(58, 8),
    to_signed(49, 8),
    to_signed(35, 8),
    to_signed(19, 8),
    to_signed(7, 8),
    to_signed(2, 8),
    to_signed(7, 8),
    to_signed(19, 8),
    to_signed(33, 8),
    to_signed(45, 8),
    to_signed(54, 8),
    to_signed(57, 8),
    to_signed(51, 8),
    to_signed(36, 8),
    to_signed(15, 8),
    to_signed(-13, 8),
    to_signed(-42, 8),
    to_signed(-70, 8),
    to_signed(-92, 8),
    to_signed(-100, 8),
    to_signed(-92, 8),
    to_signed(-70, 8),
    to_signed(-43, 8),
    to_signed(-19, 8),
    to_signed(-4, 8),
    to_signed(1, 8),
    to_signed(-4, 8),
    to_signed(-16, 8),
    to_signed(-31, 8),
    to_signed(-44, 8),
    to_signed(-49, 8),
    to_signed(-46, 8),
    to_signed(-38, 8),
    to_signed(-29, 8),
    to_signed(-18, 8),
    to_signed(-4, 8),
    to_signed(10, 8),
    to_signed(21, 8),
    to_signed(27, 8),
    to_signed(26, 8),
    to_signed(22, 8),
    to_signed(17, 8),
    to_signed(12, 8),
    to_signed(6, 8),
    to_signed(1, 8),
    to_signed(-3, 8),
    to_signed(-6, 8),
    to_signed(-11, 8),
    to_signed(-16, 8),
    to_signed(-18, 8),
    to_signed(-17, 8),
    to_signed(-14, 8),
    to_signed(-9, 8),
    to_signed(-5, 8),
    to_signed(0, 8),
    to_signed(3, 8),
    to_signed(5, 8),
    to_signed(4, 8),
    to_signed(4, 8),
    to_signed(8, 8),
    to_signed(14, 8),
    to_signed(18, 8),
    to_signed(19, 8),
    to_signed(15, 8),
    to_signed(11, 8),
    to_signed(10, 8),
    to_signed(12, 8),
    to_signed(16, 8),
    to_signed(23, 8),
    to_signed(34, 8),
    to_signed(44, 8),
    to_signed(49, 8),
    to_signed(47, 8),
    to_signed(38, 8),
    to_signed(25, 8),
    to_signed(10, 8),
    to_signed(-4, 8),
    to_signed(-14, 8),
    to_signed(-17, 8),
    to_signed(-11, 8),
    to_signed(3, 8),
    to_signed(19, 8),
    to_signed(32, 8),
    to_signed(41, 8),
    to_signed(45, 8),
    to_signed(43, 8),
    to_signed(34, 8),
    to_signed(17, 8),
    to_signed(-8, 8),
    to_signed(-37, 8),
    to_signed(-65, 8),
    to_signed(-88, 8),
    to_signed(-98, 8),
    to_signed(-88, 8),
    to_signed(-62, 8),
    to_signed(-31, 8),
    to_signed(-4, 8),
    to_signed(13, 8),
    to_signed(18, 8),
    to_signed(12, 8),
    to_signed(-3, 8),
    to_signed(-22, 8),
    to_signed(-39, 8),
    to_signed(-48, 8),
    to_signed(-45, 8),
    to_signed(-37, 8),
    to_signed(-26, 8),
    to_signed(-12, 8),
    to_signed(5, 8),
    to_signed(23, 8),
    to_signed(38, 8),
    to_signed(44, 8),
    to_signed(43, 8),
    to_signed(38, 8),
    to_signed(32, 8),
    to_signed(26, 8),
    to_signed(18, 8),
    to_signed(10, 8),
    to_signed(4, 8),
    to_signed(-2, 8),
    to_signed(-8, 8),
    to_signed(-15, 8),
    to_signed(-21, 8),
    to_signed(-23, 8),
    to_signed(-20, 8),
    to_signed(-14, 8),
    to_signed(-9, 8),
    to_signed(-6, 8),
    to_signed(-3, 8),
    to_signed(-1, 8),
    to_signed(-1, 8),
    to_signed(-3, 8),
    to_signed(-3, 8),
    to_signed(-1, 8),
    to_signed(2, 8),
    to_signed(3, 8),
    to_signed(1, 8),
    to_signed(-1, 8),
    to_signed(0, 8),
    to_signed(5, 8),
    to_signed(13, 8),
    to_signed(24, 8),
    to_signed(34, 8),
    to_signed(41, 8),
    to_signed(44, 8),
    to_signed(42, 8),
    to_signed(31, 8),
    to_signed(15, 8),
    to_signed(-2, 8),
    to_signed(-14, 8),
    to_signed(-20, 8),
    to_signed(-16, 8),
    to_signed(-3, 8),
    to_signed(17, 8),
    to_signed(36, 8),
    to_signed(52, 8),
    to_signed(61, 8),
    to_signed(63, 8),
    to_signed(59, 8),
    to_signed(48, 8),
    to_signed(33, 8),
    to_signed(11, 8),
    to_signed(-14, 8),
    to_signed(-42, 8),
    to_signed(-67, 8),
    to_signed(-81, 8),
    to_signed(-78, 8),
    to_signed(-59, 8),
    to_signed(-29, 8),
    to_signed(-1, 8),
    to_signed(17, 8),
    to_signed(24, 8),
    to_signed(20, 8),
    to_signed(8, 8),
    to_signed(-10, 8),
    to_signed(-27, 8),
    to_signed(-37, 8),
    to_signed(-38, 8),
    to_signed(-30, 8),
    to_signed(-19, 8),
    to_signed(-7, 8),
    to_signed(7, 8),
    to_signed(22, 8),
    to_signed(37, 8),
    to_signed(45, 8),
    to_signed(45, 8),
    to_signed(39, 8),
    to_signed(32, 8),
    to_signed(25, 8),
    to_signed(17, 8),
    to_signed(8, 8),
    to_signed(-1, 8),
    to_signed(-10, 8),
    to_signed(-19, 8),
    to_signed(-27, 8),
    to_signed(-34, 8),
    to_signed(-37, 8),
    to_signed(-35, 8),
    to_signed(-28, 8),
    to_signed(-19, 8),
    to_signed(-11, 8),
    to_signed(-4, 8),
    to_signed(0, 8),
    to_signed(1, 8),
    to_signed(0, 8),
    to_signed(-1, 8),
    to_signed(-2, 8),
    to_signed(-1, 8),
    to_signed(-1, 8),
    to_signed(-2, 8),
    to_signed(-2, 8),
    to_signed(-1, 8),
    to_signed(3, 8),
    to_signed(11, 8),
    to_signed(22, 8),
    to_signed(33, 8),
    to_signed(42, 8),
    to_signed(47, 8),
    to_signed(46, 8),
    to_signed(38, 8),
    to_signed(23, 8),
    to_signed(6, 8),
    to_signed(-9, 8),
    to_signed(-17, 8),
    to_signed(-14, 8),
    to_signed(-1, 8),
    to_signed(18, 8),
    to_signed(38, 8),
    to_signed(57, 8),
    to_signed(69, 8),
    to_signed(73, 8),
    to_signed(66, 8),
    to_signed(52, 8),
    to_signed(33, 8),
    to_signed(10, 8),
    to_signed(-16, 8),
    to_signed(-42, 8),
    to_signed(-65, 8),
    to_signed(-79, 8),
    to_signed(-76, 8),
    to_signed(-57, 8),
    to_signed(-30, 8),
    to_signed(-3, 8),
    to_signed(15, 8),
    to_signed(22, 8),
    to_signed(18, 8),
    to_signed(6, 8),
    to_signed(-12, 8),
    to_signed(-30, 8),
    to_signed(-43, 8),
    to_signed(-46, 8),
    to_signed(-40, 8),
    to_signed(-29, 8),
    to_signed(-16, 8),
    to_signed(-5, 8),
    to_signed(7, 8),
    to_signed(17, 8),
    to_signed(23, 8),
    to_signed(22, 8),
    to_signed(17, 8),
    to_signed(10, 8),
    to_signed(3, 8),
    to_signed(-4, 8),
    to_signed(-10, 8),
    to_signed(-16, 8),
    to_signed(-22, 8),
    to_signed(-27, 8),
    to_signed(-32, 8),
    to_signed(-36, 8),
    to_signed(-38, 8),
    to_signed(-37, 8),
    to_signed(-32, 8),
    to_signed(-26, 8),
    to_signed(-18, 8),
    to_signed(-11, 8),
    to_signed(-6, 8),
    to_signed(-3, 8),
    to_signed(-3, 8),
    to_signed(-5, 8),
    to_signed(-5, 8),
    to_signed(-4, 8),
    to_signed(-3, 8),
    to_signed(-2, 8),
    to_signed(1, 8),
    to_signed(5, 8),
    to_signed(11, 8),
    to_signed(19, 8),
    to_signed(27, 8),
    to_signed(36, 8),
    to_signed(43, 8),
    to_signed(46, 8),
    to_signed(45, 8),
    to_signed(38, 8),
    to_signed(28, 8),
    to_signed(15, 8),
    to_signed(2, 8),
    to_signed(-7, 8),
    to_signed(-8, 8),
    to_signed(1, 8),
    to_signed(17, 8),
    to_signed(33, 8),
    to_signed(45, 8),
    to_signed(55, 8),
    to_signed(59, 8),
    to_signed(56, 8),
    to_signed(46, 8),
    to_signed(30, 8),
    to_signed(10, 8),
    to_signed(-11, 8),
    to_signed(-35, 8),
    to_signed(-59, 8),
    to_signed(-78, 8),
    to_signed(-85, 8),
    to_signed(-75, 8),
    to_signed(-53, 8),
    to_signed(-29, 8),
    to_signed(-11, 8),
    to_signed(-2, 8),
    to_signed(-3, 8),
    to_signed(-11, 8),
    to_signed(-25, 8),
    to_signed(-42, 8),
    to_signed(-57, 8),
    to_signed(-65, 8),
    to_signed(-63, 8),
    to_signed(-55, 8),
    to_signed(-44, 8),
    to_signed(-31, 8),
    to_signed(-18, 8),
    to_signed(-4, 8),
    to_signed(8, 8),
    to_signed(15, 8),
    to_signed(17, 8),
    to_signed(14, 8),
    to_signed(9, 8),
    to_signed(2, 8),
    to_signed(-6, 8),
    to_signed(-14, 8),
    to_signed(-21, 8),
    to_signed(-26, 8),
    to_signed(-30, 8),
    to_signed(-33, 8),
    to_signed(-34, 8),
    to_signed(-31, 8),
    to_signed(-24, 8),
    to_signed(-14, 8),
    to_signed(-6, 8),
    to_signed(1, 8),
    to_signed(6, 8),
    to_signed(8, 8),
    to_signed(7, 8),
    to_signed(4, 8),
    to_signed(1, 8),
    to_signed(1, 8),
    to_signed(5, 8),
    to_signed(10, 8),
    to_signed(15, 8),
    to_signed(19, 8),
    to_signed(25, 8),
    to_signed(31, 8),
    to_signed(36, 8),
    to_signed(41, 8),
    to_signed(45, 8),
    to_signed(48, 8),
    to_signed(47, 8),
    to_signed(42, 8),
    to_signed(32, 8),
    to_signed(21, 8),
    to_signed(9, 8),
    to_signed(0, 8),
    to_signed(-3, 8),
    to_signed(1, 8),
    to_signed(12, 8),
    to_signed(27, 8),
    to_signed(40, 8),
    to_signed(50, 8),
    to_signed(55, 8),
    to_signed(55, 8),
    to_signed(51, 8),
    to_signed(40, 8),
    to_signed(23, 8),
    to_signed(3, 8),
    to_signed(-19, 8),
    to_signed(-44, 8),
    to_signed(-67, 8),
    to_signed(-83, 8),
    to_signed(-83, 8),
    to_signed(-68, 8),
    to_signed(-44, 8),
    to_signed(-22, 8),
    to_signed(-6, 8),
    to_signed(-1, 8),
    to_signed(-4, 8),
    to_signed(-15, 8),
    to_signed(-31, 8),
    to_signed(-48, 8),
    to_signed(-59, 8),
    to_signed(-62, 8),
    to_signed(-55, 8),
    to_signed(-44, 8),
    to_signed(-31, 8),
    to_signed(-15, 8),
    to_signed(4, 8),
    to_signed(23, 8),
    to_signed(36, 8),
    to_signed(41, 8),
    to_signed(40, 8),
    to_signed(33, 8),
    to_signed(25, 8),
    to_signed(17, 8),
    to_signed(10, 8),
    to_signed(3, 8),
    to_signed(-2, 8),
    to_signed(-5, 8),
    to_signed(-8, 8),
    to_signed(-14, 8),
    to_signed(-18, 8),
    to_signed(-16, 8),
    to_signed(-7, 8),
    to_signed(4, 8),
    to_signed(12, 8),
    to_signed(17, 8),
    to_signed(19, 8),
    to_signed(18, 8),
    to_signed(16, 8),
    to_signed(11, 8),
    to_signed(7, 8),
    to_signed(4, 8),
    to_signed(6, 8),
    to_signed(10, 8),
    to_signed(14, 8),
    to_signed(18, 8),
    to_signed(24, 8),
    to_signed(32, 8),
    to_signed(40, 8),
    to_signed(48, 8),
    to_signed(53, 8),
    to_signed(54, 8),
    to_signed(50, 8),
    to_signed(39, 8),
    to_signed(26, 8),
    to_signed(13, 8),
    to_signed(3, 8),
    to_signed(-2, 8),
    to_signed(-1, 8),
    to_signed(6, 8),
    to_signed(17, 8),
    to_signed(29, 8),
    to_signed(39, 8),
    to_signed(45, 8),
    to_signed(48, 8),
    to_signed(46, 8),
    to_signed(40, 8),
    to_signed(28, 8),
    to_signed(8, 8),
    to_signed(-15, 8),
    to_signed(-40, 8),
    to_signed(-65, 8),
    to_signed(-84, 8),
    to_signed(-93, 8),
    to_signed(-84, 8),
    to_signed(-61, 8),
    to_signed(-31, 8),
    to_signed(-5, 8),
    to_signed(11, 8),
    to_signed(14, 8),
    to_signed(5, 8),
    to_signed(-12, 8),
    to_signed(-34, 8),
    to_signed(-53, 8),
    to_signed(-65, 8),
    to_signed(-65, 8),
    to_signed(-55, 8),
    to_signed(-41, 8),
    to_signed(-24, 8),
    to_signed(-5, 8),
    to_signed(15, 8),
    to_signed(31, 8),
    to_signed(41, 8),
    to_signed(43, 8),
    to_signed(38, 8),
    to_signed(28, 8),
    to_signed(16, 8),
    to_signed(5, 8),
    to_signed(-4, 8),
    to_signed(-11, 8),
    to_signed(-15, 8),
    to_signed(-17, 8),
    to_signed(-18, 8),
    to_signed(-19, 8),
    to_signed(-17, 8),
    to_signed(-12, 8),
    to_signed(-2, 8),
    to_signed(7, 8),
    to_signed(13, 8),
    to_signed(12, 8),
    to_signed(6, 8),
    to_signed(0, 8),
    to_signed(-6, 8),
    to_signed(-9, 8),
    to_signed(-9, 8),
    to_signed(-8, 8),
    to_signed(-5, 8),
    to_signed(-1, 8),
    to_signed(4, 8),
    to_signed(11, 8),
    to_signed(19, 8),
    to_signed(29, 8),
    to_signed(39, 8),
    to_signed(48, 8),
    to_signed(54, 8),
    to_signed(52, 8),
    to_signed(42, 8),
    to_signed(25, 8),
    to_signed(5, 8),
    to_signed(-11, 8),
    to_signed(-19, 8),
    to_signed(-17, 8),
    to_signed(-7, 8),
    to_signed(7, 8),
    to_signed(24, 8),
    to_signed(40, 8),
    to_signed(51, 8),
    to_signed(54, 8),
    to_signed(49, 8),
    to_signed(40, 8),
    to_signed(27, 8),
    to_signed(11, 8),
    to_signed(-9, 8),
    to_signed(-33, 8),
    to_signed(-56, 8),
    to_signed(-76, 8),
    to_signed(-87, 8),
    to_signed(-85, 8),
    to_signed(-68, 8),
    to_signed(-41, 8),
    to_signed(-11, 8),
    to_signed(13, 8),
    to_signed(24, 8),
    to_signed(19, 8),
    to_signed(1, 8),
    to_signed(-23, 8),
    to_signed(-48, 8),
    to_signed(-64, 8),
    to_signed(-69, 8),
    to_signed(-62, 8),
    to_signed(-46, 8),
    to_signed(-24, 8),
    to_signed(1, 8),
    to_signed(25, 8),
    to_signed(44, 8),
    to_signed(54, 8),
    to_signed(55, 8),
    to_signed(48, 8),
    to_signed(35, 8),
    to_signed(20, 8),
    to_signed(6, 8),
    to_signed(-5, 8),
    to_signed(-12, 8),
    to_signed(-16, 8),
    to_signed(-18, 8),
    to_signed(-19, 8),
    to_signed(-20, 8),
    to_signed(-19, 8),
    to_signed(-15, 8),
    to_signed(-8, 8),
    to_signed(1, 8),
    to_signed(9, 8),
    to_signed(11, 8),
    to_signed(7, 8),
    to_signed(-3, 8),
    to_signed(-14, 8),
    to_signed(-21, 8),
    to_signed(-24, 8),
    to_signed(-22, 8),
    to_signed(-15, 8),
    to_signed(-6, 8),
    to_signed(3, 8),
    to_signed(10, 8),
    to_signed(16, 8),
    to_signed(22, 8),
    to_signed(27, 8),
    to_signed(31, 8),
    to_signed(34, 8),
    to_signed(35, 8),
    to_signed(30, 8),
    to_signed(18, 8),
    to_signed(3, 8),
    to_signed(-11, 8),
    to_signed(-22, 8),
    to_signed(-26, 8),
    to_signed(-20, 8),
    to_signed(-6, 8),
    to_signed(11, 8),
    to_signed(27, 8),
    to_signed(41, 8),
    to_signed(51, 8),
    to_signed(54, 8),
    to_signed(50, 8),
    to_signed(41, 8),
    to_signed(28, 8),
    to_signed(11, 8),
    to_signed(-8, 8),
    to_signed(-28, 8),
    to_signed(-47, 8),
    to_signed(-65, 8),
    to_signed(-73, 8),
    to_signed(-67, 8),
    to_signed(-48, 8),
    to_signed(-22, 8),
    to_signed(2, 8),
    to_signed(20, 8),
    to_signed(26, 8),
    to_signed(19, 8),
    to_signed(1, 8),
    to_signed(-22, 8),
    to_signed(-46, 8),
    to_signed(-62, 8),
    to_signed(-66, 8),
    to_signed(-57, 8),
    to_signed(-41, 8),
    to_signed(-20, 8),
    to_signed(6, 8),
    to_signed(33, 8),
    to_signed(53, 8),
    to_signed(61, 8),
    to_signed(56, 8),
    to_signed(43, 8),
    to_signed(24, 8),
    to_signed(7, 8),
    to_signed(-7, 8),
    to_signed(-15, 8),
    to_signed(-21, 8),
    to_signed(-25, 8),
    to_signed(-26, 8),
    to_signed(-25, 8),
    to_signed(-27, 8),
    to_signed(-26, 8),
    to_signed(-21, 8),
    to_signed(-11, 8),
    to_signed(-1, 8),
    to_signed(7, 8),
    to_signed(9, 8),
    to_signed(4, 8),
    to_signed(-7, 8),
    to_signed(-20, 8),
    to_signed(-28, 8),
    to_signed(-32, 8),
    to_signed(-31, 8),
    to_signed(-24, 8),
    to_signed(-11, 8),
    to_signed(4, 8),
    to_signed(15, 8),
    to_signed(25, 8),
    to_signed(33, 8),
    to_signed(39, 8),
    to_signed(42, 8),
    to_signed(42, 8),
    to_signed(39, 8),
    to_signed(32, 8),
    to_signed(22, 8),
    to_signed(13, 8),
    to_signed(7, 8),
    to_signed(2, 8),
    to_signed(2, 8),
    to_signed(9, 8),
    to_signed(22, 8),
    to_signed(35, 8),
    to_signed(47, 8),
    to_signed(58, 8),
    to_signed(66, 8),
    to_signed(68, 8),
    to_signed(63, 8),
    to_signed(55, 8),
    to_signed(42, 8),
    to_signed(24, 8),
    to_signed(3, 8),
    to_signed(-18, 8),
    to_signed(-37, 8),
    to_signed(-55, 8),
    to_signed(-67, 8),
    to_signed(-65, 8),
    to_signed(-52, 8),
    to_signed(-33, 8),
    to_signed(-11, 8),
    to_signed(8, 8),
    to_signed(17, 8),
    to_signed(13, 8),
    to_signed(-3, 8),
    to_signed(-25, 8),
    to_signed(-49, 8),
    to_signed(-69, 8),
    to_signed(-77, 8),
    to_signed(-71, 8),
    to_signed(-55, 8),
    to_signed(-31, 8),
    to_signed(-2, 8),
    to_signed(28, 8),
    to_signed(50, 8),
    to_signed(60, 8),
    to_signed(57, 8),
    to_signed(44, 8),
    to_signed(24, 8),
    to_signed(2, 8),
    to_signed(-15, 8),
    to_signed(-25, 8),
    to_signed(-29, 8),
    to_signed(-29, 8),
    to_signed(-27, 8),
    to_signed(-25, 8),
    to_signed(-26, 8),
    to_signed(-25, 8),
    to_signed(-19, 8),
    to_signed(-12, 8),
    to_signed(-6, 8),
    to_signed(-2, 8),
    to_signed(0, 8),
    to_signed(-3, 8),
    to_signed(-12, 8),
    to_signed(-23, 8),
    to_signed(-30, 8),
    to_signed(-30, 8),
    to_signed(-24, 8),
    to_signed(-11, 8),
    to_signed(6, 8),
    to_signed(22, 8),
    to_signed(34, 8),
    to_signed(43, 8),
    to_signed(49, 8),
    to_signed(51, 8),
    to_signed(49, 8),
    to_signed(45, 8),
    to_signed(39, 8),
    to_signed(32, 8),
    to_signed(23, 8),
    to_signed(16, 8),
    to_signed(12, 8),
    to_signed(10, 8),
    to_signed(10, 8),
    to_signed(15, 8),
    to_signed(22, 8),
    to_signed(28, 8),
    to_signed(35, 8),
    to_signed(41, 8),
    to_signed(46, 8),
    to_signed(46, 8),
    to_signed(41, 8),
    to_signed(36, 8),
    to_signed(29, 8),
    to_signed(18, 8),
    to_signed(4, 8),
    to_signed(-12, 8),
    to_signed(-30, 8),
    to_signed(-50, 8),
    to_signed(-67, 8),
    to_signed(-75, 8),
    to_signed(-72, 8),
    to_signed(-59, 8),
    to_signed(-40, 8),
    to_signed(-20, 8),
    to_signed(-7, 8),
    to_signed(-5, 8),
    to_signed(-14, 8),
    to_signed(-30, 8),
    to_signed(-51, 8),
    to_signed(-71, 8),
    to_signed(-84, 8),
    to_signed(-85, 8),
    to_signed(-74, 8),
    to_signed(-55, 8),
    to_signed(-29, 8),
    to_signed(0, 8),
    to_signed(26, 8),
    to_signed(44, 8),
    to_signed(51, 8),
    to_signed(48, 8),
    to_signed(36, 8),
    to_signed(19, 8),
    to_signed(3, 8),
    to_signed(-7, 8),
    to_signed(-10, 8),
    to_signed(-10, 8),
    to_signed(-9, 8),
    to_signed(-8, 8),
    to_signed(-6, 8),
    to_signed(-4, 8),
    to_signed(2, 8),
    to_signed(10, 8),
    to_signed(17, 8),
    to_signed(20, 8),
    to_signed(18, 8),
    to_signed(11, 8),
    to_signed(-1, 8),
    to_signed(-15, 8),
    to_signed(-26, 8),
    to_signed(-29, 8),
    to_signed(-24, 8),
    to_signed(-13, 8),
    to_signed(4, 8),
    to_signed(21, 8),
    to_signed(34, 8),
    to_signed(42, 8),
    to_signed(45, 8),
    to_signed(45, 8),
    to_signed(42, 8),
    to_signed(36, 8),
    to_signed(29, 8),
    to_signed(24, 8),
    to_signed(20, 8),
    to_signed(18, 8),
    to_signed(18, 8),
    to_signed(17, 8),
    to_signed(13, 8),
    to_signed(8, 8),
    to_signed(5, 8),
    to_signed(6, 8),
    to_signed(10, 8),
    to_signed(16, 8),
    to_signed(26, 8),
    to_signed(36, 8),
    to_signed(41, 8),
    to_signed(41, 8),
    to_signed(35, 8),
    to_signed(23, 8),
    to_signed(5, 8),
    to_signed(-17, 8),
    to_signed(-41, 8),
    to_signed(-67, 8),
    to_signed(-89, 8),
    to_signed(-102, 8),
    to_signed(-96, 8),
    to_signed(-73, 8),
    to_signed(-42, 8),
    to_signed(-14, 8),
    to_signed(6, 8),
    to_signed(13, 8),
    to_signed(6, 8),
    to_signed(-11, 8),
    to_signed(-35, 8),
    to_signed(-60, 8),
    to_signed(-78, 8),
    to_signed(-81, 8),
    to_signed(-69, 8),
    to_signed(-45, 8),
    to_signed(-16, 8),
    to_signed(16, 8),
    to_signed(47, 8),
    to_signed(71, 8),
    to_signed(79, 8),
    to_signed(72, 8),
    to_signed(55, 8),
    to_signed(32, 8),
    to_signed(10, 8),
    to_signed(-5, 8),
    to_signed(-10, 8),
    to_signed(-11, 8),
    to_signed(-10, 8),
    to_signed(-8, 8),
    to_signed(-5, 8),
    to_signed(-3, 8),
    to_signed(-1, 8),
    to_signed(4, 8),
    to_signed(11, 8),
    to_signed(14, 8),
    to_signed(10, 8),
    to_signed(1, 8),
    to_signed(-12, 8),
    to_signed(-29, 8),
    to_signed(-44, 8),
    to_signed(-51, 8),
    to_signed(-49, 8),
    to_signed(-39, 8),
    to_signed(-23, 8),
    to_signed(-2, 8),
    to_signed(20, 8),
    to_signed(35, 8),
    to_signed(41, 8),
    to_signed(42, 8),
    to_signed(38, 8),
    to_signed(29, 8),
    to_signed(18, 8),
    to_signed(10, 8),
    to_signed(5, 8),
    to_signed(2, 8),
    to_signed(0, 8),
    to_signed(0, 8),
    to_signed(-2, 8),
    to_signed(-6, 8),
    to_signed(-7, 8),
    to_signed(-1, 8),
    to_signed(10, 8),
    to_signed(23, 8),
    to_signed(37, 8),
    to_signed(51, 8),
    to_signed(59, 8),
    to_signed(58, 8),
    to_signed(50, 8),
    to_signed(37, 8),
    to_signed(20, 8),
    to_signed(-2, 8),
    to_signed(-24, 8),
    to_signed(-45, 8),
    to_signed(-65, 8),
    to_signed(-77, 8),
    to_signed(-72, 8),
    to_signed(-50, 8),
    to_signed(-21, 8),
    to_signed(5, 8),
    to_signed(21, 8),
    to_signed(24, 8),
    to_signed(14, 8),
    to_signed(-6, 8),
    to_signed(-29, 8),
    to_signed(-52, 8),
    to_signed(-69, 8),
    to_signed(-73, 8),
    to_signed(-61, 8),
    to_signed(-38, 8),
    to_signed(-10, 8),
    to_signed(21, 8),
    to_signed(50, 8),
    to_signed(73, 8),
    to_signed(81, 8),
    to_signed(74, 8),
    to_signed(57, 8),
    to_signed(33, 8),
    to_signed(9, 8),
    to_signed(-8, 8),
    to_signed(-15, 8),
    to_signed(-17, 8),
    to_signed(-18, 8),
    to_signed(-18, 8),
    to_signed(-18, 8),
    to_signed(-18, 8),
    to_signed(-18, 8),
    to_signed(-14, 8),
    to_signed(-7, 8),
    to_signed(-2, 8),
    to_signed(-2, 8),
    to_signed(-7, 8),
    to_signed(-18, 8),
    to_signed(-32, 8),
    to_signed(-47, 8),
    to_signed(-55, 8),
    to_signed(-56, 8),
    to_signed(-50, 8),
    to_signed(-36, 8),
    to_signed(-14, 8),
    to_signed(12, 8),
    to_signed(35, 8),
    to_signed(51, 8),
    to_signed(58, 8),
    to_signed(56, 8),
    to_signed(45, 8),
    to_signed(32, 8),
    to_signed(20, 8),
    to_signed(13, 8),
    to_signed(9, 8),
    to_signed(8, 8),
    to_signed(10, 8),
    to_signed(10, 8),
    to_signed(10, 8),
    to_signed(13, 8),
    to_signed(21, 8),
    to_signed(32, 8),
    to_signed(43, 8),
    to_signed(53, 8),
    to_signed(62, 8),
    to_signed(65, 8),
    to_signed(60, 8),
    to_signed(50, 8),
    to_signed(36, 8),
    to_signed(20, 8),
    to_signed(4, 8),
    to_signed(-11, 8),
    to_signed(-26, 8),
    to_signed(-42, 8),
    to_signed(-55, 8),
    to_signed(-59, 8),
    to_signed(-49, 8),
    to_signed(-32, 8),
    to_signed(-14, 8),
    to_signed(-2, 8),
    to_signed(3, 8),
    to_signed(-2, 8),
    to_signed(-15, 8),
    to_signed(-31, 8),
    to_signed(-48, 8),
    to_signed(-61, 8),
    to_signed(-65, 8),
    to_signed(-56, 8),
    to_signed(-40, 8),
    to_signed(-21, 8),
    to_signed(-1, 8),
    to_signed(21, 8),
    to_signed(40, 8),
    to_signed(50, 8),
    to_signed(49, 8),
    to_signed(39, 8),
    to_signed(23, 8),
    to_signed(7, 8),
    to_signed(-7, 8),
    to_signed(-16, 8),
    to_signed(-22, 8),
    to_signed(-25, 8),
    to_signed(-25, 8),
    to_signed(-24, 8),
    to_signed(-24, 8),
    to_signed(-26, 8),
    to_signed(-23, 8),
    to_signed(-14, 8),
    to_signed(-6, 8),
    to_signed(-5, 8),
    to_signed(-9, 8),
    to_signed(-17, 8),
    to_signed(-28, 8),
    to_signed(-39, 8),
    to_signed(-45, 8),
    to_signed(-44, 8),
    to_signed(-39, 8),
    to_signed(-26, 8),
    to_signed(-6, 8),
    to_signed(17, 8),
    to_signed(37, 8),
    to_signed(49, 8),
    to_signed(55, 8),
    to_signed(55, 8),
    to_signed(48, 8),
    to_signed(36, 8),
    to_signed(25, 8),
    to_signed(19, 8),
    to_signed(16, 8),
    to_signed(16, 8),
    to_signed(18, 8),
    to_signed(17, 8),
    to_signed(14, 8),
    to_signed(11, 8),
    to_signed(13, 8),
    to_signed(17, 8),
    to_signed(21, 8),
    to_signed(27, 8),
    to_signed(35, 8),
    to_signed(43, 8),
    to_signed(46, 8),
    to_signed(43, 8),
    to_signed(34, 8),
    to_signed(22, 8),
    to_signed(10, 8),
    to_signed(0, 8),
    to_signed(-10, 8),
    to_signed(-24, 8),
    to_signed(-42, 8),
    to_signed(-57, 8),
    to_signed(-63, 8),
    to_signed(-58, 8),
    to_signed(-47, 8),
    to_signed(-34, 8),
    to_signed(-22, 8),
    to_signed(-14, 8),
    to_signed(-14, 8),
    to_signed(-22, 8),
    to_signed(-36, 8),
    to_signed(-52, 8),
    to_signed(-63, 8),
    to_signed(-66, 8),
    to_signed(-61, 8),
    to_signed(-50, 8),
    to_signed(-37, 8),
    to_signed(-18, 8),
    to_signed(5, 8),
    to_signed(26, 8),
    to_signed(40, 8),
    to_signed(45, 8),
    to_signed(44, 8),
    to_signed(38, 8),
    to_signed(28, 8),
    to_signed(16, 8),
    to_signed(4, 8),
    to_signed(-7, 8),
    to_signed(-14, 8),
    to_signed(-18, 8),
    to_signed(-20, 8),
    to_signed(-21, 8),
    to_signed(-20, 8),
    to_signed(-15, 8),
    to_signed(-5, 8),
    to_signed(5, 8),
    to_signed(8, 8),
    to_signed(4, 8),
    to_signed(-6, 8),
    to_signed(-19, 8),
    to_signed(-30, 8),
    to_signed(-36, 8),
    to_signed(-35, 8),
    to_signed(-27, 8),
    to_signed(-12, 8),
    to_signed(9, 8),
    to_signed(33, 8),
    to_signed(51, 8),
    to_signed(60, 8),
    to_signed(62, 8),
    to_signed(59, 8),
    to_signed(51, 8),
    to_signed(41, 8),
    to_signed(33, 8),
    to_signed(27, 8),
    to_signed(24, 8),
    to_signed(22, 8),
    to_signed(19, 8),
    to_signed(13, 8),
    to_signed(4, 8),
    to_signed(-2, 8),
    to_signed(-2, 8),
    to_signed(4, 8),
    to_signed(13, 8),
    to_signed(25, 8),
    to_signed(37, 8),
    to_signed(48, 8),
    to_signed(52, 8),
    to_signed(48, 8),
    to_signed(37, 8),
    to_signed(21, 8),
    to_signed(4, 8),
    to_signed(-11, 8),
    to_signed(-27, 8),
    to_signed(-46, 8),
    to_signed(-66, 8),
    to_signed(-77, 8),
    to_signed(-73, 8),
    to_signed(-55, 8),
    to_signed(-30, 8),
    to_signed(-8, 8),
    to_signed(7, 8),
    to_signed(11, 8),
    to_signed(5, 8),
    to_signed(-9, 8),
    to_signed(-29, 8),
    to_signed(-47, 8),
    to_signed(-58, 8),
    to_signed(-57, 8),
    to_signed(-47, 8),
    to_signed(-33, 8),
    to_signed(-14, 8),
    to_signed(9, 8),
    to_signed(34, 8),
    to_signed(55, 8),
    to_signed(64, 8),
    to_signed(63, 8),
    to_signed(56, 8),
    to_signed(45, 8),
    to_signed(32, 8),
    to_signed(19, 8),
    to_signed(6, 8),
    to_signed(-5, 8),
    to_signed(-11, 8),
    to_signed(-12, 8),
    to_signed(-12, 8),
    to_signed(-12, 8),
    to_signed(-12, 8),
    to_signed(-8, 8),
    to_signed(-2, 8),
    to_signed(6, 8),
    to_signed(9, 8),
    to_signed(4, 8),
    to_signed(-7, 8),
    to_signed(-20, 8),
    to_signed(-31, 8),
    to_signed(-37, 8),
    to_signed(-38, 8),
    to_signed(-31, 8),
    to_signed(-17, 8),
    to_signed(2, 8),
    to_signed(22, 8),
    to_signed(36, 8),
    to_signed(41, 8),
    to_signed(40, 8),
    to_signed(37, 8),
    to_signed(33, 8),
    to_signed(28, 8),
    to_signed(24, 8),
    to_signed(21, 8),
    to_signed(18, 8),
    to_signed(15, 8),
    to_signed(10, 8),
    to_signed(4, 8),
    to_signed(-2, 8),
    to_signed(-1, 8),
    to_signed(6, 8),
    to_signed(17, 8),
    to_signed(28, 8),
    to_signed(36, 8),
    to_signed(43, 8),
    to_signed(46, 8),
    to_signed(44, 8),
    to_signed(38, 8),
    to_signed(28, 8),
    to_signed(15, 8),
    to_signed(1, 8),
    to_signed(-14, 8),
    to_signed(-34, 8),
    to_signed(-59, 8),
    to_signed(-79, 8),
    to_signed(-85, 8),
    to_signed(-71, 8),
    to_signed(-45, 8),
    to_signed(-17, 8),
    to_signed(5, 8),
    to_signed(17, 8),
    to_signed(16, 8),
    to_signed(3, 8),
    to_signed(-16, 8),
    to_signed(-39, 8),
    to_signed(-57, 8),
    to_signed(-65, 8),
    to_signed(-61, 8),
    to_signed(-50, 8),
    to_signed(-34, 8),
    to_signed(-11, 8),
    to_signed(17, 8),
    to_signed(42, 8),
    to_signed(58, 8),
    to_signed(63, 8),
    to_signed(60, 8),
    to_signed(49, 8),
    to_signed(35, 8),
    to_signed(20, 8),
    to_signed(6, 8),
    to_signed(-8, 8),
    to_signed(-19, 8),
    to_signed(-24, 8),
    to_signed(-24, 8),
    to_signed(-24, 8),
    to_signed(-23, 8),
    to_signed(-21, 8),
    to_signed(-16, 8),
    to_signed(-10, 8),
    to_signed(-5, 8),
    to_signed(-3, 8),
    to_signed(-7, 8),
    to_signed(-17, 8),
    to_signed(-30, 8),
    to_signed(-39, 8),
    to_signed(-43, 8),
    to_signed(-41, 8),
    to_signed(-31, 8),
    to_signed(-13, 8),
    to_signed(9, 8),
    to_signed(27, 8),
    to_signed(38, 8),
    to_signed(42, 8),
    to_signed(41, 8),
    to_signed(38, 8),
    to_signed(35, 8),
    to_signed(30, 8),
    to_signed(22, 8),
    to_signed(12, 8),
    to_signed(4, 8),
    to_signed(-2, 8),
    to_signed(-5, 8),
    to_signed(-6, 8),
    to_signed(-3, 8),
    to_signed(6, 8),
    to_signed(18, 8),
    to_signed(28, 8),
    to_signed(35, 8),
    to_signed(39, 8),
    to_signed(42, 8),
    to_signed(42, 8),
    to_signed(39, 8),
    to_signed(32, 8),
    to_signed(21, 8),
    to_signed(9, 8),
    to_signed(-3, 8),
    to_signed(-17, 8),
    to_signed(-38, 8),
    to_signed(-62, 8),
    to_signed(-79, 8),
    to_signed(-79, 8),
    to_signed(-65, 8),
    to_signed(-42, 8),
    to_signed(-19, 8),
    to_signed(-1, 8),
    to_signed(8, 8),
    to_signed(4, 8),
    to_signed(-12, 8),
    to_signed(-34, 8),
    to_signed(-56, 8),
    to_signed(-70, 8),
    to_signed(-71, 8),
    to_signed(-61, 8),
    to_signed(-44, 8),
    to_signed(-23, 8),
    to_signed(3, 8),
    to_signed(30, 8),
    to_signed(48, 8),
    to_signed(56, 8),
    to_signed(55, 8),
    to_signed(49, 8),
    to_signed(39, 8),
    to_signed(25, 8),
    to_signed(9, 8),
    to_signed(-8, 8),
    to_signed(-23, 8),
    to_signed(-33, 8),
    to_signed(-36, 8),
    to_signed(-35, 8),
    to_signed(-33, 8),
    to_signed(-30, 8),
    to_signed(-23, 8),
    to_signed(-15, 8),
    to_signed(-8, 8),
    to_signed(-4, 8),
    to_signed(-4, 8),
    to_signed(-9, 8),
    to_signed(-20, 8),
    to_signed(-30, 8),
    to_signed(-36, 8),
    to_signed(-35, 8),
    to_signed(-28, 8),
    to_signed(-13, 8),
    to_signed(7, 8),
    to_signed(26, 8),
    to_signed(37, 8),
    to_signed(40, 8),
    to_signed(37, 8),
    to_signed(33, 8),
    to_signed(31, 8),
    to_signed(31, 8),
    to_signed(29, 8),
    to_signed(24, 8),
    to_signed(17, 8),
    to_signed(10, 8),
    to_signed(3, 8),
    to_signed(-3, 8),
    to_signed(-9, 8),
    to_signed(-10, 8),
    to_signed(-6, 8),
    to_signed(2, 8),
    to_signed(13, 8),
    to_signed(25, 8),
    to_signed(37, 8),
    to_signed(48, 8),
    to_signed(54, 8),
    to_signed(51, 8),
    to_signed(40, 8),
    to_signed(24, 8),
    to_signed(8, 8),
    to_signed(-6, 8),
    to_signed(-23, 8),
    to_signed(-46, 8),
    to_signed(-69, 8),
    to_signed(-84, 8),
    to_signed(-82, 8),
    to_signed(-64, 8),
    to_signed(-37, 8),
    to_signed(-9, 8),
    to_signed(13, 8),
    to_signed(24, 8),
    to_signed(19, 8),
    to_signed(-3, 8),
    to_signed(-31, 8),
    to_signed(-55, 8),
    to_signed(-66, 8),
    to_signed(-66, 8),
    to_signed(-55, 8),
    to_signed(-37, 8),
    to_signed(-12, 8),
    to_signed(16, 8),
    to_signed(41, 8),
    to_signed(56, 8),
    to_signed(61, 8),
    to_signed(59, 8),
    to_signed(53, 8),
    to_signed(43, 8),
    to_signed(28, 8),
    to_signed(10, 8),
    to_signed(-8, 8),
    to_signed(-23, 8),
    to_signed(-32, 8),
    to_signed(-35, 8),
    to_signed(-33, 8),
    to_signed(-26, 8),
    to_signed(-18, 8),
    to_signed(-8, 8),
    to_signed(1, 8),
    to_signed(7, 8),
    to_signed(8, 8),
    to_signed(2, 8),
    to_signed(-8, 8),
    to_signed(-22, 8),
    to_signed(-34, 8),
    to_signed(-39, 8),
    to_signed(-34, 8),
    to_signed(-21, 8),
    to_signed(-2, 8),
    to_signed(20, 8),
    to_signed(39, 8),
    to_signed(51, 8),
    to_signed(54, 8),
    to_signed(50, 8),
    to_signed(43, 8),
    to_signed(37, 8),
    to_signed(33, 8),
    to_signed(31, 8),
    to_signed(27, 8),
    to_signed(23, 8),
    to_signed(19, 8),
    to_signed(16, 8),
    to_signed(12, 8),
    to_signed(6, 8),
    to_signed(2, 8),
    to_signed(4, 8),
    to_signed(10, 8),
    to_signed(21, 8),
    to_signed(34, 8),
    to_signed(48, 8),
    to_signed(59, 8),
    to_signed(66, 8),
    to_signed(64, 8),
    to_signed(53, 8),
    to_signed(37, 8),
    to_signed(21, 8),
    to_signed(5, 8),
    to_signed(-14, 8),
    to_signed(-37, 8),
    to_signed(-57, 8),
    to_signed(-65, 8),
    to_signed(-58, 8),
    to_signed(-40, 8),
    to_signed(-16, 8),
    to_signed(7, 8),
    to_signed(23, 8),
    to_signed(26, 8),
    to_signed(15, 8),
    to_signed(-9, 8),
    to_signed(-36, 8),
    to_signed(-56, 8),
    to_signed(-63, 8),
    to_signed(-60, 8),
    to_signed(-49, 8),
    to_signed(-31, 8),
    to_signed(-5, 8),
    to_signed(23, 8),
    to_signed(46, 8),
    to_signed(59, 8),
    to_signed(62, 8),
    to_signed(57, 8),
    to_signed(46, 8),
    to_signed(33, 8),
    to_signed(18, 8),
    to_signed(2, 8),
    to_signed(-13, 8),
    to_signed(-23, 8),
    to_signed(-30, 8),
    to_signed(-32, 8),
    to_signed(-32, 8),
    to_signed(-27, 8),
    to_signed(-19, 8),
    to_signed(-12, 8),
    to_signed(-8, 8),
    to_signed(-6, 8),
    to_signed(-6, 8),
    to_signed(-10, 8),
    to_signed(-19, 8),
    to_signed(-30, 8),
    to_signed(-38, 8),
    to_signed(-39, 8),
    to_signed(-32, 8),
    to_signed(-16, 8),
    to_signed(6, 8),
    to_signed(31, 8),
    to_signed(50, 8),
    to_signed(61, 8),
    to_signed(61, 8),
    to_signed(53, 8),
    to_signed(42, 8),
    to_signed(33, 8),
    to_signed(29, 8),
    to_signed(26, 8),
    to_signed(24, 8),
    to_signed(21, 8),
    to_signed(18, 8),
    to_signed(14, 8),
    to_signed(7, 8),
    to_signed(1, 8),
    to_signed(-2, 8),
    to_signed(0, 8),
    to_signed(8, 8),
    to_signed(20, 8),
    to_signed(33, 8),
    to_signed(45, 8),
    to_signed(53, 8),
    to_signed(56, 8),
    to_signed(54, 8),
    to_signed(42, 8),
    to_signed(27, 8),
    to_signed(11, 8),
    to_signed(-6, 8),
    to_signed(-28, 8),
    to_signed(-52, 8),
    to_signed(-69, 8),
    to_signed(-73, 8),
    to_signed(-63, 8),
    to_signed(-45, 8),
    to_signed(-24, 8),
    to_signed(-6, 8),
    to_signed(4, 8),
    to_signed(5, 8),
    to_signed(-6, 8),
    to_signed(-28, 8),
    to_signed(-55, 8),
    to_signed(-74, 8),
    to_signed(-80, 8),
    to_signed(-74, 8),
    to_signed(-62, 8),
    to_signed(-41, 8),
    to_signed(-11, 8),
    to_signed(19, 8),
    to_signed(41, 8),
    to_signed(53, 8),
    to_signed(54, 8),
    to_signed(47, 8),
    to_signed(35, 8),
    to_signed(21, 8),
    to_signed(6, 8),
    to_signed(-10, 8),
    to_signed(-24, 8),
    to_signed(-33, 8),
    to_signed(-37, 8),
    to_signed(-38, 8),
    to_signed(-36, 8),
    to_signed(-27, 8),
    to_signed(-15, 8),
    to_signed(-4, 8),
    to_signed(3, 8),
    to_signed(6, 8),
    to_signed(3, 8),
    to_signed(-6, 8),
    to_signed(-17, 8),
    to_signed(-28, 8),
    to_signed(-35, 8),
    to_signed(-36, 8),
    to_signed(-27, 8),
    to_signed(-10, 8),
    to_signed(12, 8),
    to_signed(31, 8),
    to_signed(44, 8),
    to_signed(50, 8),
    to_signed(49, 8),
    to_signed(41, 8),
    to_signed(33, 8),
    to_signed(26, 8),
    to_signed(24, 8),
    to_signed(23, 8),
    to_signed(22, 8),
    to_signed(19, 8),
    to_signed(14, 8),
    to_signed(7, 8),
    to_signed(0, 8),
    to_signed(-4, 8),
    to_signed(-5, 8),
    to_signed(-3, 8),
    to_signed(5, 8),
    to_signed(18, 8),
    to_signed(32, 8),
    to_signed(43, 8),
    to_signed(47, 8),
    to_signed(44, 8),
    to_signed(33, 8),
    to_signed(17, 8),
    to_signed(-1, 8),
    to_signed(-18, 8),
    to_signed(-37, 8),
    to_signed(-57, 8),
    to_signed(-76, 8),
    to_signed(-86, 8),
    to_signed(-82, 8),
    to_signed(-66, 8),
    to_signed(-43, 8),
    to_signed(-20, 8),
    to_signed(-5, 8),
    to_signed(2, 8),
    to_signed(-1, 8),
    to_signed(-14, 8),
    to_signed(-34, 8),
    to_signed(-54, 8),
    to_signed(-67, 8),
    to_signed(-69, 8),
    to_signed(-61, 8),
    to_signed(-46, 8),
    to_signed(-25, 8),
    to_signed(0, 8),
    to_signed(25, 8),
    to_signed(43, 8),
    to_signed(52, 8),
    to_signed(54, 8),
    to_signed(50, 8),
    to_signed(41, 8),
    to_signed(28, 8),
    to_signed(13, 8),
    to_signed(-2, 8),
    to_signed(-16, 8),
    to_signed(-25, 8),
    to_signed(-31, 8),
    to_signed(-33, 8),
    to_signed(-32, 8),
    to_signed(-26, 8),
    to_signed(-15, 8),
    to_signed(-2, 8),
    to_signed(8, 8),
    to_signed(11, 8),
    to_signed(6, 8),
    to_signed(-6, 8),
    to_signed(-22, 8),
    to_signed(-35, 8),
    to_signed(-42, 8),
    to_signed(-44, 8),
    to_signed(-36, 8),
    to_signed(-20, 8),
    to_signed(0, 8),
    to_signed(17, 8),
    to_signed(28, 8),
    to_signed(32, 8),
    to_signed(31, 8),
    to_signed(27, 8),
    to_signed(23, 8),
    to_signed(21, 8),
    to_signed(21, 8),
    to_signed(21, 8),
    to_signed(21, 8),
    to_signed(17, 8),
    to_signed(10, 8),
    to_signed(1, 8),
    to_signed(-7, 8),
    to_signed(-12, 8),
    to_signed(-12, 8),
    to_signed(-6, 8),
    to_signed(8, 8),
    to_signed(28, 8),
    to_signed(48, 8),
    to_signed(63, 8),
    to_signed(66, 8),
    to_signed(57, 8),
    to_signed(43, 8),
    to_signed(28, 8),
    to_signed(14, 8),
    to_signed(0, 8),
    to_signed(-13, 8),
    to_signed(-29, 8),
    to_signed(-46, 8),
    to_signed(-58, 8),
    to_signed(-58, 8),
    to_signed(-45, 8),
    to_signed(-24, 8),
    to_signed(-4, 8),
    to_signed(9, 8),
    to_signed(13, 8),
    to_signed(7, 8),
    to_signed(-8, 8),
    to_signed(-27, 8),
    to_signed(-47, 8),
    to_signed(-61, 8),
    to_signed(-65, 8),
    to_signed(-57, 8),
    to_signed(-41, 8),
    to_signed(-22, 8),
    to_signed(1, 8),
    to_signed(25, 8),
    to_signed(45, 8),
    to_signed(54, 8),
    to_signed(55, 8),
    to_signed(49, 8),
    to_signed(38, 8),
    to_signed(23, 8),
    to_signed(7, 8),
    to_signed(-8, 8),
    to_signed(-20, 8),
    to_signed(-29, 8),
    to_signed(-33, 8),
    to_signed(-33, 8),
    to_signed(-32, 8),
    to_signed(-28, 8),
    to_signed(-19, 8),
    to_signed(-7, 8),
    to_signed(2, 8),
    to_signed(5, 8),
    to_signed(0, 8),
    to_signed(-10, 8),
    to_signed(-22, 8),
    to_signed(-31, 8),
    to_signed(-34, 8),
    to_signed(-30, 8),
    to_signed(-21, 8),
    to_signed(-3, 8),
    to_signed(19, 8),
    to_signed(37, 8),
    to_signed(43, 8),
    to_signed(42, 8),
    to_signed(38, 8),
    to_signed(33, 8),
    to_signed(29, 8),
    to_signed(26, 8),
    to_signed(25, 8),
    to_signed(25, 8),
    to_signed(23, 8),
    to_signed(20, 8),
    to_signed(16, 8),
    to_signed(9, 8),
    to_signed(1, 8),
    to_signed(-5, 8),
    to_signed(-8, 8),
    to_signed(-4, 8),
    to_signed(8, 8),
    to_signed(28, 8),
    to_signed(48, 8),
    to_signed(60, 8),
    to_signed(63, 8),
    to_signed(58, 8),
    to_signed(47, 8),
    to_signed(32, 8),
    to_signed(17, 8),
    to_signed(5, 8),
    to_signed(-6, 8),
    to_signed(-20, 8),
    to_signed(-38, 8),
    to_signed(-53, 8),
    to_signed(-59, 8),
    to_signed(-52, 8),
    to_signed(-35, 8),
    to_signed(-17, 8),
    to_signed(-2, 8),
    to_signed(5, 8),
    to_signed(3, 8),
    to_signed(-8, 8),
    to_signed(-26, 8),
    to_signed(-46, 8),
    to_signed(-59, 8),
    to_signed(-62, 8),
    to_signed(-57, 8),
    to_signed(-45, 8),
    to_signed(-28, 8),
    to_signed(-6, 8),
    to_signed(18, 8),
    to_signed(38, 8),
    to_signed(50, 8),
    to_signed(55, 8),
    to_signed(51, 8),
    to_signed(43, 8),
    to_signed(30, 8),
    to_signed(16, 8),
    to_signed(1, 8),
    to_signed(-14, 8),
    to_signed(-26, 8),
    to_signed(-31, 8),
    to_signed(-33, 8),
    to_signed(-34, 8),
    to_signed(-32, 8),
    to_signed(-26, 8),
    to_signed(-15, 8),
    to_signed(-4, 8),
    to_signed(2, 8),
    to_signed(1, 8),
    to_signed(-8, 8),
    to_signed(-21, 8),
    to_signed(-34, 8),
    to_signed(-41, 8),
    to_signed(-42, 8),
    to_signed(-34, 8),
    to_signed(-16, 8),
    to_signed(5, 8),
    to_signed(23, 8),
    to_signed(30, 8),
    to_signed(29, 8),
    to_signed(25, 8),
    to_signed(22, 8),
    to_signed(23, 8),
    to_signed(27, 8),
    to_signed(30, 8),
    to_signed(29, 8),
    to_signed(24, 8),
    to_signed(16, 8),
    to_signed(6, 8),
    to_signed(-4, 8),
    to_signed(-14, 8),
    to_signed(-20, 8),
    to_signed(-18, 8),
    to_signed(-8, 8),
    to_signed(9, 8),
    to_signed(29, 8),
    to_signed(46, 8),
    to_signed(56, 8),
    to_signed(58, 8),
    to_signed(55, 8),
    to_signed(45, 8),
    to_signed(31, 8),
    to_signed(19, 8),
    to_signed(11, 8),
    to_signed(5, 8),
    to_signed(-8, 8),
    to_signed(-28, 8),
    to_signed(-48, 8),
    to_signed(-58, 8),
    to_signed(-52, 8),
    to_signed(-33, 8),
    to_signed(-10, 8),
    to_signed(9, 8),
    to_signed(19, 8),
    to_signed(19, 8),
    to_signed(7, 8),
    to_signed(-17, 8),
    to_signed(-44, 8),
    to_signed(-63, 8),
    to_signed(-70, 8),
    to_signed(-68, 8),
    to_signed(-60, 8),
    to_signed(-45, 8),
    to_signed(-21, 8),
    to_signed(5, 8),
    to_signed(28, 8),
    to_signed(42, 8),
    to_signed(48, 8),
    to_signed(48, 8),
    to_signed(41, 8),
    to_signed(26, 8),
    to_signed(5, 8),
    to_signed(-16, 8),
    to_signed(-31, 8),
    to_signed(-40, 8),
    to_signed(-44, 8),
    to_signed(-44, 8),
    to_signed(-42, 8),
    to_signed(-38, 8),
    to_signed(-31, 8),
    to_signed(-20, 8),
    to_signed(-9, 8),
    to_signed(-1, 8),
    to_signed(0, 8),
    to_signed(-6, 8),
    to_signed(-19, 8),
    to_signed(-33, 8),
    to_signed(-44, 8),
    to_signed(-49, 8),
    to_signed(-45, 8),
    to_signed(-30, 8),
    to_signed(-6, 8),
    to_signed(18, 8),
    to_signed(34, 8),
    to_signed(42, 8),
    to_signed(44, 8),
    to_signed(43, 8),
    to_signed(43, 8),
    to_signed(45, 8),
    to_signed(48, 8),
    to_signed(46, 8),
    to_signed(39, 8),
    to_signed(30, 8),
    to_signed(23, 8),
    to_signed(17, 8),
    to_signed(10, 8),
    to_signed(5, 8),
    to_signed(5, 8),
    to_signed(14, 8),
    to_signed(31, 8),
    to_signed(51, 8),
    to_signed(68, 8),
    to_signed(78, 8),
    to_signed(82, 8),
    to_signed(80, 8),
    to_signed(69, 8),
    to_signed(51, 8),
    to_signed(33, 8),
    to_signed(22, 8),
    to_signed(12, 8),
    to_signed(-4, 8),
    to_signed(-28, 8),
    to_signed(-50, 8),
    to_signed(-62, 8),
    to_signed(-60, 8),
    to_signed(-47, 8),
    to_signed(-26, 8),
    to_signed(-5, 8),
    to_signed(10, 8),
    to_signed(14, 8),
    to_signed(4, 8),
    to_signed(-19, 8),
    to_signed(-47, 8),
    to_signed(-71, 8),
    to_signed(-85, 8),
    to_signed(-89, 8),
    to_signed(-85, 8),
    to_signed(-70, 8),
    to_signed(-44, 8),
    to_signed(-13, 8),
    to_signed(17, 8),
    to_signed(39, 8),
    to_signed(53, 8),
    to_signed(56, 8),
    to_signed(48, 8),
    to_signed(29, 8),
    to_signed(4, 8),
    to_signed(-21, 8),
    to_signed(-40, 8),
    to_signed(-48, 8),
    to_signed(-46, 8),
    to_signed(-39, 8),
    to_signed(-28, 8),
    to_signed(-15, 8),
    to_signed(-1, 8),
    to_signed(10, 8),
    to_signed(15, 8),
    to_signed(16, 8),
    to_signed(14, 8),
    to_signed(7, 8),
    to_signed(-5, 8),
    to_signed(-19, 8),
    to_signed(-28, 8),
    to_signed(-29, 8),
    to_signed(-25, 8),
    to_signed(-14, 8),
    to_signed(2, 8),
    to_signed(22, 8),
    to_signed(39, 8),
    to_signed(49, 8),
    to_signed(52, 8),
    to_signed(52, 8),
    to_signed(54, 8),
    to_signed(57, 8),
    to_signed(54, 8),
    to_signed(45, 8),
    to_signed(31, 8),
    to_signed(20, 8),
    to_signed(12, 8),
    to_signed(4, 8),
    to_signed(-4, 8),
    to_signed(-8, 8),
    to_signed(-6, 8),
    to_signed(5, 8),
    to_signed(19, 8),
    to_signed(35, 8),
    to_signed(48, 8),
    to_signed(57, 8),
    to_signed(62, 8),
    to_signed(61, 8),
    to_signed(53, 8),
    to_signed(39, 8),
    to_signed(24, 8),
    to_signed(11, 8),
    to_signed(0, 8),
    to_signed(-15, 8),
    to_signed(-35, 8),
    to_signed(-56, 8),
    to_signed(-70, 8),
    to_signed(-70, 8),
    to_signed(-57, 8),
    to_signed(-37, 8),
    to_signed(-15, 8),
    to_signed(2, 8),
    to_signed(10, 8),
    to_signed(4, 8),
    to_signed(-15, 8),
    to_signed(-39, 8),
    to_signed(-59, 8),
    to_signed(-72, 8),
    to_signed(-79, 8),
    to_signed(-77, 8),
    to_signed(-64, 8),
    to_signed(-38, 8),
    to_signed(-5, 8),
    to_signed(28, 8),
    to_signed(55, 8),
    to_signed(72, 8),
    to_signed(78, 8),
    to_signed(72, 8),
    to_signed(54, 8),
    to_signed(28, 8),
    to_signed(3, 8),
    to_signed(-17, 8),
    to_signed(-28, 8),
    to_signed(-32, 8),
    to_signed(-26, 8),
    to_signed(-15, 8),
    to_signed(-4, 8),
    to_signed(3, 8),
    to_signed(6, 8),
    to_signed(9, 8),
    to_signed(11, 8),
    to_signed(10, 8),
    to_signed(4, 8),
    to_signed(-4, 8),
    to_signed(-13, 8),
    to_signed(-20, 8),
    to_signed(-23, 8),
    to_signed(-21, 8),
    to_signed(-15, 8),
    to_signed(-5, 8),
    to_signed(11, 8),
    to_signed(28, 8),
    to_signed(41, 8),
    to_signed(47, 8),
    to_signed(50, 8),
    to_signed(50, 8),
    to_signed(47, 8),
    to_signed(41, 8),
    to_signed(33, 8),
    to_signed(22, 8),
    to_signed(11, 8),
    to_signed(1, 8),
    to_signed(-9, 8),
    to_signed(-20, 8),
    to_signed(-28, 8),
    to_signed(-28, 8),
    to_signed(-17, 8),
    to_signed(1, 8),
    to_signed(19, 8),
    to_signed(36, 8),
    to_signed(49, 8),
    to_signed(58, 8),
    to_signed(57, 8),
    to_signed(48, 8),
    to_signed(33, 8),
    to_signed(21, 8),
    to_signed(15, 8),
    to_signed(10, 8),
    to_signed(2, 8),
    to_signed(-12, 8),
    to_signed(-30, 8),
    to_signed(-49, 8),
    to_signed(-62, 8),
    to_signed(-63, 8),
    to_signed(-50, 8),
    to_signed(-29, 8),
    to_signed(-7, 8),
    to_signed(8, 8),
    to_signed(12, 8),
    to_signed(4, 8),
    to_signed(-14, 8),
    to_signed(-37, 8),
    to_signed(-60, 8),
    to_signed(-77, 8),
    to_signed(-83, 8),
    to_signed(-76, 8),
    to_signed(-56, 8),
    to_signed(-26, 8),
    to_signed(9, 8),
    to_signed(42, 8),
    to_signed(66, 8),
    to_signed(74, 8),
    to_signed(69, 8),
    to_signed(53, 8),
    to_signed(30, 8),
    to_signed(3, 8),
    to_signed(-18, 8),
    to_signed(-29, 8),
    to_signed(-33, 8),
    to_signed(-29, 8),
    to_signed(-20, 8),
    to_signed(-9, 8),
    to_signed(-4, 8),
    to_signed(-5, 8),
    to_signed(-7, 8),
    to_signed(-8, 8),
    to_signed(-11, 8),
    to_signed(-16, 8),
    to_signed(-22, 8),
    to_signed(-27, 8),
    to_signed(-33, 8),
    to_signed(-36, 8),
    to_signed(-37, 8),
    to_signed(-34, 8),
    to_signed(-28, 8),
    to_signed(-15, 8),
    to_signed(3, 8),
    to_signed(18, 8),
    to_signed(27, 8),
    to_signed(32, 8),
    to_signed(35, 8),
    to_signed(35, 8),
    to_signed(29, 8),
    to_signed(23, 8),
    to_signed(19, 8),
    to_signed(15, 8),
    to_signed(9, 8),
    to_signed(4, 8),
    to_signed(0, 8),
    to_signed(-4, 8),
    to_signed(-8, 8),
    to_signed(-8, 8),
    to_signed(-2, 8),
    to_signed(8, 8),
    to_signed(20, 8),
    to_signed(34, 8),
    to_signed(47, 8),
    to_signed(54, 8),
    to_signed(56, 8),
    to_signed(53, 8),
    to_signed(47, 8),
    to_signed(37, 8),
    to_signed(29, 8),
    to_signed(20, 8),
    to_signed(9, 8),
    to_signed(-9, 8),
    to_signed(-29, 8),
    to_signed(-47, 8),
    to_signed(-56, 8),
    to_signed(-53, 8),
    to_signed(-36, 8),
    to_signed(-12, 8),
    to_signed(10, 8),
    to_signed(23, 8),
    to_signed(23, 8),
    to_signed(11, 8),
    to_signed(-11, 8),
    to_signed(-38, 8),
    to_signed(-62, 8),
    to_signed(-77, 8),
    to_signed(-78, 8),
    to_signed(-68, 8),
    to_signed(-48, 8),
    to_signed(-22, 8),
    to_signed(11, 8),
    to_signed(41, 8),
    to_signed(58, 8),
    to_signed(59, 8),
    to_signed(48, 8),
    to_signed(34, 8),
    to_signed(16, 8),
    to_signed(-3, 8),
    to_signed(-21, 8),
    to_signed(-33, 8),
    to_signed(-37, 8),
    to_signed(-36, 8),
    to_signed(-34, 8),
    to_signed(-33, 8),
    to_signed(-33, 8),
    to_signed(-29, 8),
    to_signed(-22, 8),
    to_signed(-17, 8),
    to_signed(-15, 8),
    to_signed(-16, 8),
    to_signed(-20, 8),
    to_signed(-30, 8),
    to_signed(-41, 8),
    to_signed(-49, 8),
    to_signed(-48, 8),
    to_signed(-42, 8),
    to_signed(-32, 8),
    to_signed(-16, 8),
    to_signed(3, 8),
    to_signed(19, 8),
    to_signed(29, 8),
    to_signed(37, 8),
    to_signed(43, 8),
    to_signed(45, 8),
    to_signed(41, 8),
    to_signed(35, 8),
    to_signed(26, 8),
    to_signed(17, 8),
    to_signed(7, 8),
    to_signed(1, 8),
    to_signed(-4, 8),
    to_signed(-9, 8),
    to_signed(-10, 8),
    to_signed(-4, 8),
    to_signed(8, 8),
    to_signed(20, 8),
    to_signed(35, 8),
    to_signed(50, 8),
    to_signed(61, 8),
    to_signed(64, 8),
    to_signed(61, 8),
    to_signed(53, 8),
    to_signed(41, 8),
    to_signed(25, 8),
    to_signed(12, 8),
    to_signed(1, 8),
    to_signed(-13, 8),
    to_signed(-34, 8),
    to_signed(-56, 8),
    to_signed(-67, 8),
    to_signed(-63, 8),
    to_signed(-45, 8),
    to_signed(-20, 8),
    to_signed(5, 8),
    to_signed(21, 8),
    to_signed(23, 8),
    to_signed(8, 8),
    to_signed(-19, 8),
    to_signed(-51, 8),
    to_signed(-77, 8),
    to_signed(-89, 8),
    to_signed(-86, 8),
    to_signed(-73, 8),
    to_signed(-53, 8),
    to_signed(-24, 8),
    to_signed(9, 8),
    to_signed(37, 8),
    to_signed(54, 8),
    to_signed(56, 8),
    to_signed(46, 8),
    to_signed(30, 8),
    to_signed(12, 8),
    to_signed(-6, 8),
    to_signed(-22, 8),
    to_signed(-34, 8),
    to_signed(-38, 8),
    to_signed(-33, 8),
    to_signed(-25, 8),
    to_signed(-19, 8),
    to_signed(-15, 8),
    to_signed(-10, 8),
    to_signed(-4, 8),
    to_signed(0, 8),
    to_signed(1, 8),
    to_signed(-1, 8),
    to_signed(-6, 8),
    to_signed(-13, 8),
    to_signed(-22, 8),
    to_signed(-30, 8),
    to_signed(-32, 8),
    to_signed(-28, 8),
    to_signed(-18, 8),
    to_signed(-2, 8),
    to_signed(19, 8),
    to_signed(40, 8),
    to_signed(56, 8),
    to_signed(65, 8),
    to_signed(67, 8),
    to_signed(62, 8),
    to_signed(53, 8),
    to_signed(41, 8),
    to_signed(28, 8),
    to_signed(15, 8),
    to_signed(7, 8),
    to_signed(4, 8),
    to_signed(3, 8),
    to_signed(1, 8),
    to_signed(1, 8),
    to_signed(4, 8),
    to_signed(12, 8),
    to_signed(21, 8),
    to_signed(28, 8),
    to_signed(35, 8),
    to_signed(40, 8),
    to_signed(41, 8),
    to_signed(36, 8),
    to_signed(26, 8),
    to_signed(17, 8),
    to_signed(8, 8),
    to_signed(2, 8),
    to_signed(-3, 8),
    to_signed(-8, 8),
    to_signed(-19, 8),
    to_signed(-36, 8),
    to_signed(-54, 8),
    to_signed(-64, 8),
    to_signed(-62, 8),
    to_signed(-50, 8),
    to_signed(-30, 8),
    to_signed(-10, 8),
    to_signed(4, 8),
    to_signed(7, 8),
    to_signed(-3, 8),
    to_signed(-25, 8),
    to_signed(-49, 8),
    to_signed(-68, 8),
    to_signed(-74, 8),
    to_signed(-70, 8),
    to_signed(-56, 8),
    to_signed(-34, 8),
    to_signed(-4, 8),
    to_signed(28, 8),
    to_signed(52, 8),
    to_signed(63, 8),
    to_signed(62, 8),
    to_signed(53, 8),
    to_signed(38, 8),
    to_signed(19, 8),
    to_signed(1, 8),
    to_signed(-13, 8),
    to_signed(-19, 8),
    to_signed(-19, 8),
    to_signed(-13, 8),
    to_signed(-5, 8),
    to_signed(1, 8),
    to_signed(2, 8),
    to_signed(0, 8),
    to_signed(-2, 8),
    to_signed(-5, 8),
    to_signed(-7, 8),
    to_signed(-11, 8),
    to_signed(-17, 8),
    to_signed(-25, 8),
    to_signed(-34, 8),
    to_signed(-41, 8),
    to_signed(-42, 8),
    to_signed(-37, 8),
    to_signed(-23, 8),
    to_signed(-2, 8),
    to_signed(19, 8),
    to_signed(34, 8),
    to_signed(43, 8),
    to_signed(45, 8),
    to_signed(41, 8),
    to_signed(32, 8),
    to_signed(23, 8),
    to_signed(15, 8),
    to_signed(8, 8),
    to_signed(2, 8),
    to_signed(-1, 8),
    to_signed(-1, 8),
    to_signed(0, 8),
    to_signed(0, 8),
    to_signed(2, 8),
    to_signed(6, 8),
    to_signed(13, 8),
    to_signed(21, 8),
    to_signed(31, 8),
    to_signed(40, 8),
    to_signed(48, 8),
    to_signed(52, 8),
    to_signed(52, 8),
    to_signed(46, 8),
    to_signed(36, 8),
    to_signed(25, 8),
    to_signed(17, 8),
    to_signed(9, 8),
    to_signed(0, 8),
    to_signed(-13, 8),
    to_signed(-27, 8),
    to_signed(-39, 8),
    to_signed(-46, 8),
    to_signed(-44, 8),
    to_signed(-35, 8),
    to_signed(-21, 8),
    to_signed(-8, 8),
    to_signed(0, 8),
    to_signed(0, 8),
    to_signed(-9, 8),
    to_signed(-27, 8),
    to_signed(-46, 8),
    to_signed(-60, 8),
    to_signed(-64, 8),
    to_signed(-58, 8),
    to_signed(-44, 8),
    to_signed(-24, 8),
    to_signed(2, 8),
    to_signed(27, 8),
    to_signed(46, 8),
    to_signed(53, 8),
    to_signed(52, 8),
    to_signed(45, 8),
    to_signed(34, 8),
    to_signed(20, 8),
    to_signed(4, 8),
    to_signed(-9, 8),
    to_signed(-17, 8),
    to_signed(-19, 8),
    to_signed(-20, 8),
    to_signed(-20, 8),
    to_signed(-22, 8),
    to_signed(-24, 8),
    to_signed(-24, 8),
    to_signed(-19, 8),
    to_signed(-13, 8),
    to_signed(-8, 8),
    to_signed(-8, 8),
    to_signed(-13, 8),
    to_signed(-22, 8),
    to_signed(-31, 8),
    to_signed(-36, 8),
    to_signed(-36, 8),
    to_signed(-29, 8),
    to_signed(-13, 8),
    to_signed(9, 8),
    to_signed(30, 8),
    to_signed(45, 8),
    to_signed(53, 8),
    to_signed(58, 8),
    to_signed(57, 8),
    to_signed(51, 8),
    to_signed(42, 8),
    to_signed(32, 8),
    to_signed(24, 8),
    to_signed(16, 8),
    to_signed(10, 8),
    to_signed(7, 8),
    to_signed(5, 8),
    to_signed(4, 8),
    to_signed(5, 8),
    to_signed(7, 8),
    to_signed(11, 8),
    to_signed(18, 8),
    to_signed(27, 8),
    to_signed(35, 8),
    to_signed(40, 8),
    to_signed(43, 8),
    to_signed(42, 8),
    to_signed(35, 8),
    to_signed(24, 8),
    to_signed(13, 8),
    to_signed(4, 8),
    to_signed(-4, 8),
    to_signed(-15, 8),
    to_signed(-28, 8),
    to_signed(-39, 8),
    to_signed(-46, 8),
    to_signed(-48, 8),
    to_signed(-44, 8),
    to_signed(-34, 8),
    to_signed(-19, 8),
    to_signed(-5, 8),
    to_signed(1, 8),
    to_signed(-4, 8),
    to_signed(-21, 8),
    to_signed(-41, 8),
    to_signed(-60, 8),
    to_signed(-71, 8),
    to_signed(-72, 8),
    to_signed(-61, 8),
    to_signed(-41, 8),
    to_signed(-16, 8),
    to_signed(10, 8),
    to_signed(32, 8),
    to_signed(45, 8),
    to_signed(49, 8),
    to_signed(47, 8),
    to_signed(41, 8),
    to_signed(31, 8),
    to_signed(18, 8),
    to_signed(2, 8),
    to_signed(-10, 8),
    to_signed(-17, 8),
    to_signed(-18, 8),
    to_signed(-16, 8),
    to_signed(-14, 8),
    to_signed(-13, 8),
    to_signed(-10, 8),
    to_signed(-6, 8),
    to_signed(-4, 8),
    to_signed(-6, 8),
    to_signed(-10, 8),
    to_signed(-15, 8),
    to_signed(-20, 8),
    to_signed(-27, 8),
    to_signed(-31, 8),
    to_signed(-28, 8),
    to_signed(-19, 8),
    to_signed(-6, 8),
    to_signed(7, 8),
    to_signed(21, 8),
    to_signed(33, 8),
    to_signed(41, 8),
    to_signed(47, 8),
    to_signed(51, 8),
    to_signed(51, 8),
    to_signed(48, 8),
    to_signed(42, 8),
    to_signed(34, 8),
    to_signed(25, 8),
    to_signed(18, 8),
    to_signed(12, 8),
    to_signed(7, 8),
    to_signed(2, 8),
    to_signed(-1, 8),
    to_signed(0, 8),
    to_signed(2, 8),
    to_signed(5, 8),
    to_signed(10, 8),
    to_signed(16, 8),
    to_signed(23, 8),
    to_signed(26, 8),
    to_signed(26, 8),
    to_signed(23, 8),
    to_signed(19, 8),
    to_signed(15, 8),
    to_signed(14, 8),
    to_signed(14, 8),
    to_signed(15, 8),
    to_signed(12, 8),
    to_signed(4, 8),
    to_signed(-9, 8),
    to_signed(-26, 8),
    to_signed(-41, 8),
    to_signed(-49, 8),
    to_signed(-46, 8),
    to_signed(-34, 8),
    to_signed(-18, 8),
    to_signed(-7, 8),
    to_signed(-3, 8),
    to_signed(-7, 8),
    to_signed(-14, 8),
    to_signed(-25, 8),
    to_signed(-37, 8),
    to_signed(-47, 8),
    to_signed(-49, 8),
    to_signed(-43, 8),
    to_signed(-29, 8),
    to_signed(-13, 8),
    to_signed(5, 8),
    to_signed(24, 8),
    to_signed(40, 8),
    to_signed(50, 8),
    to_signed(52, 8),
    to_signed(44, 8),
    to_signed(31, 8),
    to_signed(15, 8),
    to_signed(1, 8),
    to_signed(-8, 8),
    to_signed(-13, 8),
    to_signed(-12, 8),
    to_signed(-10, 8),
    to_signed(-9, 8),
    to_signed(-9, 8),
    to_signed(-9, 8),
    to_signed(-11, 8),
    to_signed(-16, 8),
    to_signed(-21, 8),
    to_signed(-25, 8),
    to_signed(-28, 8),
    to_signed(-30, 8),
    to_signed(-29, 8),
    to_signed(-25, 8),
    to_signed(-20, 8),
    to_signed(-14, 8),
    to_signed(-8, 8),
    to_signed(-1, 8),
    to_signed(8, 8),
    to_signed(18, 8),
    to_signed(27, 8),
    to_signed(32, 8),
    to_signed(33, 8),
    to_signed(30, 8),
    to_signed(25, 8),
    to_signed(22, 8),
    to_signed(19, 8),
    to_signed(18, 8),
    to_signed(15, 8),
    to_signed(11, 8),
    to_signed(4, 8),
    to_signed(-2, 8),
    to_signed(-7, 8),
    to_signed(-10, 8),
    to_signed(-10, 8),
    to_signed(-5, 8),
    to_signed(7, 8),
    to_signed(21, 8),
    to_signed(33, 8),
    to_signed(40, 8),
    to_signed(43, 8),
    to_signed(44, 8),
    to_signed(43, 8),
    to_signed(39, 8),
    to_signed(33, 8),
    to_signed(28, 8),
    to_signed(22, 8),
    to_signed(9, 8),
    to_signed(-13, 8),
    to_signed(-39, 8),
    to_signed(-58, 8),
    to_signed(-64, 8),
    to_signed(-57, 8),
    to_signed(-40, 8),
    to_signed(-21, 8),
    to_signed(-3, 8),
    to_signed(9, 8),
    to_signed(13, 8),
    to_signed(5, 8),
    to_signed(-13, 8),
    to_signed(-35, 8),
    to_signed(-51, 8),
    to_signed(-58, 8),
    to_signed(-55, 8),
    to_signed(-44, 8),
    to_signed(-26, 8),
    to_signed(-4, 8),
    to_signed(17, 8),
    to_signed(35, 8),
    to_signed(46, 8),
    to_signed(49, 8),
    to_signed(45, 8),
    to_signed(37, 8),
    to_signed(26, 8),
    to_signed(14, 8),
    to_signed(2, 8),
    to_signed(-8, 8),
    to_signed(-16, 8),
    to_signed(-25, 8),
    to_signed(-34, 8),
    to_signed(-42, 8),
    to_signed(-46, 8),
    to_signed(-46, 8),
    to_signed(-42, 8),
    to_signed(-36, 8),
    to_signed(-30, 8),
    to_signed(-23, 8),
    to_signed(-20, 8),
    to_signed(-20, 8),
    to_signed(-23, 8),
    to_signed(-28, 8),
    to_signed(-29, 8),
    to_signed(-26, 8),
    to_signed(-18, 8),
    to_signed(-6, 8),
    to_signed(8, 8),
    to_signed(20, 8),
    to_signed(28, 8),
    to_signed(30, 8),
    to_signed(30, 8),
    to_signed(31, 8),
    to_signed(33, 8),
    to_signed(32, 8),
    to_signed(27, 8),
    to_signed(21, 8),
    to_signed(14, 8),
    to_signed(6, 8),
    to_signed(-3, 8),
    to_signed(-12, 8),
    to_signed(-16, 8),
    to_signed(-12, 8),
    to_signed(2, 8),
    to_signed(22, 8),
    to_signed(45, 8),
    to_signed(64, 8),
    to_signed(76, 8),
    to_signed(80, 8),
    to_signed(75, 8),
    to_signed(59, 8),
    to_signed(40, 8),
    to_signed(23, 8),
    to_signed(8, 8),
    to_signed(-9, 8),
    to_signed(-31, 8),
    to_signed(-57, 8),
    to_signed(-75, 8),
    to_signed(-78, 8),
    to_signed(-64, 8),
    to_signed(-40, 8),
    to_signed(-14, 8),
    to_signed(5, 8),
    to_signed(15, 8),
    to_signed(12, 8),
    to_signed(-5, 8),
    to_signed(-32, 8),
    to_signed(-57, 8),
    to_signed(-72, 8),
    to_signed(-72, 8),
    to_signed(-61, 8),
    to_signed(-43, 8),
    to_signed(-20, 8),
    to_signed(4, 8),
    to_signed(26, 8),
    to_signed(40, 8),
    to_signed(47, 8),
    to_signed(45, 8),
    to_signed(39, 8),
    to_signed(30, 8),
    to_signed(19, 8),
    to_signed(7, 8),
    to_signed(-5, 8),
    to_signed(-14, 8),
    to_signed(-22, 8),
    to_signed(-31, 8),
    to_signed(-42, 8),
    to_signed(-51, 8),
    to_signed(-55, 8),
    to_signed(-54, 8),
    to_signed(-46, 8),
    to_signed(-36, 8),
    to_signed(-26, 8),
    to_signed(-18, 8),
    to_signed(-14, 8),
    to_signed(-13, 8),
    to_signed(-16, 8),
    to_signed(-18, 8),
    to_signed(-17, 8),
    to_signed(-13, 8),
    to_signed(-4, 8),
    to_signed(8, 8),
    to_signed(20, 8),
    to_signed(32, 8),
    to_signed(39, 8),
    to_signed(43, 8),
    to_signed(44, 8),
    to_signed(44, 8),
    to_signed(42, 8),
    to_signed(37, 8),
    to_signed(30, 8),
    to_signed(21, 8),
    to_signed(13, 8),
    to_signed(8, 8),
    to_signed(3, 8),
    to_signed(-3, 8),
    to_signed(-6, 8),
    to_signed(-2, 8),
    to_signed(10, 8),
    to_signed(28, 8),
    to_signed(46, 8),
    to_signed(61, 8),
    to_signed(70, 8),
    to_signed(71, 8),
    to_signed(63, 8),
    to_signed(49, 8),
    to_signed(33, 8),
    to_signed(22, 8),
    to_signed(16, 8),
    to_signed(7, 8),
    to_signed(-12, 8),
    to_signed(-38, 8),
    to_signed(-60, 8),
    to_signed(-68, 8),
    to_signed(-61, 8),
    to_signed(-42, 8),
    to_signed(-20, 8),
    to_signed(-2, 8),
    to_signed(4, 8),
    to_signed(-1, 8),
    to_signed(-16, 8),
    to_signed(-37, 8),
    to_signed(-58, 8),
    to_signed(-70, 8),
    to_signed(-70, 8),
    to_signed(-61, 8),
    to_signed(-47, 8),
    to_signed(-28, 8),
    to_signed(-7, 8),
    to_signed(13, 8),
    to_signed(29, 8),
    to_signed(39, 8),
    to_signed(41, 8),
    to_signed(38, 8),
    to_signed(33, 8),
    to_signed(28, 8),
    to_signed(20, 8),
    to_signed(10, 8),
    to_signed(-1, 8),
    to_signed(-11, 8),
    to_signed(-21, 8),
    to_signed(-32, 8),
    to_signed(-41, 8),
    to_signed(-45, 8),
    to_signed(-42, 8),
    to_signed(-35, 8),
    to_signed(-26, 8),
    to_signed(-19, 8),
    to_signed(-15, 8),
    to_signed(-15, 8),
    to_signed(-17, 8),
    to_signed(-19, 8),
    to_signed(-21, 8),
    to_signed(-17, 8),
    to_signed(-8, 8),
    to_signed(4, 8),
    to_signed(18, 8),
    to_signed(32, 8),
    to_signed(44, 8),
    to_signed(50, 8),
    to_signed(51, 8),
    to_signed(47, 8),
    to_signed(41, 8),
    to_signed(35, 8),
    to_signed(27, 8),
    to_signed(21, 8),
    to_signed(16, 8),
    to_signed(13, 8),
    to_signed(11, 8),
    to_signed(7, 8),
    to_signed(0, 8),
    to_signed(-7, 8),
    to_signed(-10, 8),
    to_signed(-6, 8),
    to_signed(4, 8),
    to_signed(17, 8),
    to_signed(30, 8),
    to_signed(42, 8),
    to_signed(49, 8),
    to_signed(49, 8),
    to_signed(45, 8),
    to_signed(39, 8),
    to_signed(32, 8),
    to_signed(26, 8),
    to_signed(16, 8),
    to_signed(-2, 8),
    to_signed(-29, 8),
    to_signed(-57, 8),
    to_signed(-76, 8),
    to_signed(-77, 8),
    to_signed(-63, 8),
    to_signed(-41, 8),
    to_signed(-21, 8),
    to_signed(-8, 8),
    to_signed(-4, 8),
    to_signed(-10, 8),
    to_signed(-23, 8),
    to_signed(-40, 8),
    to_signed(-56, 8),
    to_signed(-64, 8),
    to_signed(-61, 8),
    to_signed(-51, 8),
    to_signed(-36, 8),
    to_signed(-16, 8),
    to_signed(8, 8),
    to_signed(30, 8),
    to_signed(46, 8),
    to_signed(55, 8),
    to_signed(56, 8),
    to_signed(53, 8),
    to_signed(46, 8),
    to_signed(36, 8),
    to_signed(25, 8),
    to_signed(12, 8),
    to_signed(0, 8),
    to_signed(-10, 8),
    to_signed(-19, 8),
    to_signed(-26, 8),
    to_signed(-30, 8),
    to_signed(-28, 8),
    to_signed(-22, 8),
    to_signed(-12, 8),
    to_signed(-3, 8),
    to_signed(2, 8),
    to_signed(2, 8),
    to_signed(-4, 8),
    to_signed(-11, 8),
    to_signed(-17, 8),
    to_signed(-20, 8),
    to_signed(-17, 8),
    to_signed(-9, 8),
    to_signed(1, 8),
    to_signed(13, 8),
    to_signed(25, 8),
    to_signed(34, 8),
    to_signed(38, 8),
    to_signed(38, 8),
    to_signed(34, 8),
    to_signed(30, 8),
    to_signed(26, 8),
    to_signed(22, 8),
    to_signed(16, 8),
    to_signed(10, 8),
    to_signed(5, 8),
    to_signed(0, 8),
    to_signed(-5, 8),
    to_signed(-8, 8),
    to_signed(-8, 8),
    to_signed(-2, 8),
    to_signed(11, 8),
    to_signed(27, 8),
    to_signed(42, 8),
    to_signed(52, 8),
    to_signed(57, 8),
    to_signed(56, 8),
    to_signed(50, 8),
    to_signed(41, 8),
    to_signed(32, 8),
    to_signed(24, 8),
    to_signed(16, 8),
    to_signed(3, 8),
    to_signed(-18, 8),
    to_signed(-44, 8),
    to_signed(-67, 8),
    to_signed(-75, 8),
    to_signed(-64, 8),
    to_signed(-40, 8),
    to_signed(-12, 8),
    to_signed(9, 8),
    to_signed(19, 8),
    to_signed(18, 8),
    to_signed(7, 8),
    to_signed(-12, 8),
    to_signed(-35, 8),
    to_signed(-52, 8),
    to_signed(-59, 8),
    to_signed(-54, 8),
    to_signed(-42, 8),
    to_signed(-23, 8),
    to_signed(0, 8),
    to_signed(24, 8),
    to_signed(45, 8),
    to_signed(58, 8),
    to_signed(63, 8),
    to_signed(59, 8),
    to_signed(51, 8),
    to_signed(41, 8),
    to_signed(29, 8),
    to_signed(15, 8),
    to_signed(2, 8),
    to_signed(-9, 8),
    to_signed(-17, 8),
    to_signed(-25, 8),
    to_signed(-29, 8),
    to_signed(-28, 8),
    to_signed(-21, 8),
    to_signed(-12, 8),
    to_signed(-4, 8),
    to_signed(-1, 8),
    to_signed(-5, 8),
    to_signed(-16, 8),
    to_signed(-29, 8),
    to_signed(-40, 8),
    to_signed(-43, 8),
    to_signed(-37, 8),
    to_signed(-24, 8),
    to_signed(-7, 8),
    to_signed(9, 8),
    to_signed(24, 8),
    to_signed(37, 8),
    to_signed(44, 8),
    to_signed(45, 8),
    to_signed(44, 8),
    to_signed(41, 8),
    to_signed(37, 8),
    to_signed(32, 8),
    to_signed(28, 8),
    to_signed(22, 8),
    to_signed(14, 8),
    to_signed(7, 8),
    to_signed(-1, 8),
    to_signed(-7, 8),
    to_signed(-11, 8),
    to_signed(-8, 8),
    to_signed(2, 8),
    to_signed(19, 8),
    to_signed(37, 8),
    to_signed(50, 8),
    to_signed(56, 8),
    to_signed(54, 8),
    to_signed(47, 8),
    to_signed(38, 8),
    to_signed(30, 8),
    to_signed(21, 8),
    to_signed(14, 8),
    to_signed(4, 8),
    to_signed(-13, 8),
    to_signed(-37, 8),
    to_signed(-61, 8),
    to_signed(-75, 8),
    to_signed(-72, 8),
    to_signed(-54, 8),
    to_signed(-31, 8),
    to_signed(-9, 8),
    to_signed(3, 8),
    to_signed(5, 8),
    to_signed(-3, 8),
    to_signed(-21, 8),
    to_signed(-43, 8),
    to_signed(-62, 8),
    to_signed(-71, 8),
    to_signed(-67, 8),
    to_signed(-54, 8),
    to_signed(-35, 8),
    to_signed(-10, 8),
    to_signed(18, 8),
    to_signed(43, 8),
    to_signed(59, 8),
    to_signed(64, 8),
    to_signed(59, 8),
    to_signed(47, 8),
    to_signed(31, 8),
    to_signed(15, 8),
    to_signed(0, 8),
    to_signed(-12, 8),
    to_signed(-19, 8),
    to_signed(-24, 8),
    to_signed(-29, 8),
    to_signed(-36, 8),
    to_signed(-39, 8),
    to_signed(-36, 8),
    to_signed(-29, 8),
    to_signed(-21, 8),
    to_signed(-16, 8),
    to_signed(-15, 8),
    to_signed(-18, 8),
    to_signed(-24, 8),
    to_signed(-30, 8),
    to_signed(-33, 8),
    to_signed(-31, 8),
    to_signed(-23, 8),
    to_signed(-12, 8),
    to_signed(0, 8),
    to_signed(10, 8),
    to_signed(19, 8),
    to_signed(27, 8),
    to_signed(31, 8),
    to_signed(30, 8),
    to_signed(26, 8),
    to_signed(21, 8),
    to_signed(16, 8),
    to_signed(11, 8),
    to_signed(7, 8),
    to_signed(3, 8),
    to_signed(-2, 8),
    to_signed(-7, 8),
    to_signed(-10, 8),
    to_signed(-8, 8),
    to_signed(0, 8),
    to_signed(13, 8),
    to_signed(30, 8),
    to_signed(48, 8),
    to_signed(60, 8),
    to_signed(65, 8),
    to_signed(63, 8),
    to_signed(54, 8),
    to_signed(42, 8),
    to_signed(32, 8),
    to_signed(25, 8),
    to_signed(20, 8),
    to_signed(13, 8),
    to_signed(-1, 8),
    to_signed(-23, 8),
    to_signed(-51, 8),
    to_signed(-73, 8),
    to_signed(-81, 8),
    to_signed(-73, 8),
    to_signed(-55, 8),
    to_signed(-34, 8),
    to_signed(-15, 8),
    to_signed(-4, 8),
    to_signed(-4, 8),
    to_signed(-15, 8),
    to_signed(-32, 8),
    to_signed(-51, 8),
    to_signed(-65, 8),
    to_signed(-71, 8),
    to_signed(-68, 8),
    to_signed(-57, 8),
    to_signed(-38, 8),
    to_signed(-11, 8),
    to_signed(18, 8),
    to_signed(38, 8),
    to_signed(47, 8),
    to_signed(46, 8),
    to_signed(39, 8),
    to_signed(26, 8),
    to_signed(10, 8),
    to_signed(-4, 8),
    to_signed(-14, 8),
    to_signed(-20, 8),
    to_signed(-23, 8),
    to_signed(-25, 8),
    to_signed(-29, 8),
    to_signed(-34, 8),
    to_signed(-34, 8),
    to_signed(-28, 8),
    to_signed(-22, 8),
    to_signed(-20, 8),
    to_signed(-19, 8),
    to_signed(-19, 8),
    to_signed(-23, 8),
    to_signed(-30, 8),
    to_signed(-36, 8),
    to_signed(-37, 8),
    to_signed(-33, 8),
    to_signed(-22, 8),
    to_signed(-6, 8),
    to_signed(9, 8),
    to_signed(21, 8),
    to_signed(30, 8),
    to_signed(36, 8),
    to_signed(39, 8),
    to_signed(36, 8),
    to_signed(32, 8),
    to_signed(28, 8),
    to_signed(26, 8),
    to_signed(24, 8),
    to_signed(21, 8),
    to_signed(18, 8),
    to_signed(11, 8),
    to_signed(3, 8),
    to_signed(-3, 8),
    to_signed(-4, 8),
    to_signed(1, 8),
    to_signed(11, 8),
    to_signed(25, 8),
    to_signed(37, 8),
    to_signed(45, 8),
    to_signed(46, 8),
    to_signed(42, 8),
    to_signed(34, 8),
    to_signed(25, 8),
    to_signed(18, 8),
    to_signed(16, 8),
    to_signed(14, 8),
    to_signed(4, 8),
    to_signed(-17, 8),
    to_signed(-44, 8),
    to_signed(-70, 8),
    to_signed(-87, 8),
    to_signed(-89, 8),
    to_signed(-77, 8),
    to_signed(-57, 8),
    to_signed(-37, 8),
    to_signed(-21, 8),
    to_signed(-14, 8),
    to_signed(-21, 8),
    to_signed(-37, 8),
    to_signed(-56, 8),
    to_signed(-70, 8),
    to_signed(-78, 8),
    to_signed(-77, 8),
    to_signed(-67, 8),
    to_signed(-48, 8),
    to_signed(-21, 8),
    to_signed(10, 8),
    to_signed(37, 8),
    to_signed(55, 8),
    to_signed(62, 8),
    to_signed(62, 8),
    to_signed(55, 8),
    to_signed(43, 8),
    to_signed(29, 8),
    to_signed(17, 8),
    to_signed(9, 8),
    to_signed(2, 8),
    to_signed(-6, 8),
    to_signed(-15, 8),
    to_signed(-24, 8),
    to_signed(-28, 8),
    to_signed(-26, 8),
    to_signed(-20, 8),
    to_signed(-14, 8),
    to_signed(-10, 8),
    to_signed(-6, 8),
    to_signed(-3, 8),
    to_signed(-5, 8),
    to_signed(-11, 8),
    to_signed(-15, 8),
    to_signed(-15, 8),
    to_signed(-11, 8),
    to_signed(-3, 8),
    to_signed(8, 8),
    to_signed(20, 8),
    to_signed(29, 8),
    to_signed(35, 8),
    to_signed(39, 8),
    to_signed(40, 8),
    to_signed(36, 8),
    to_signed(30, 8),
    to_signed(24, 8),
    to_signed(18, 8),
    to_signed(11, 8),
    to_signed(5, 8),
    to_signed(-1, 8),
    to_signed(-8, 8),
    to_signed(-14, 8),
    to_signed(-17, 8),
    to_signed(-12, 8),
    to_signed(-1, 8),
    to_signed(14, 8),
    to_signed(32, 8),
    to_signed(48, 8),
    to_signed(60, 8),
    to_signed(64, 8),
    to_signed(61, 8),
    to_signed(52, 8),
    to_signed(38, 8),
    to_signed(23, 8),
    to_signed(9, 8),
    to_signed(-6, 8),
    to_signed(-29, 8),
    to_signed(-56, 8),
    to_signed(-79, 8),
    to_signed(-88, 8),
    to_signed(-81, 8),
    to_signed(-59, 8),
    to_signed(-31, 8),
    to_signed(-6, 8),
    to_signed(8, 8),
    to_signed(9, 8),
    to_signed(-2, 8),
    to_signed(-24, 8),
    to_signed(-48, 8),
    to_signed(-65, 8),
    to_signed(-69, 8),
    to_signed(-62, 8),
    to_signed(-48, 8),
    to_signed(-26, 8),
    to_signed(4, 8),
    to_signed(35, 8),
    to_signed(60, 8),
    to_signed(75, 8),
    to_signed(79, 8),
    to_signed(72, 8),
    to_signed(58, 8),
    to_signed(41, 8),
    to_signed(25, 8),
    to_signed(13, 8),
    to_signed(5, 8),
    to_signed(1, 8),
    to_signed(-3, 8),
    to_signed(-8, 8),
    to_signed(-13, 8),
    to_signed(-14, 8),
    to_signed(-12, 8),
    to_signed(-10, 8),
    to_signed(-9, 8),
    to_signed(-8, 8),
    to_signed(-7, 8),
    to_signed(-7, 8),
    to_signed(-12, 8),
    to_signed(-20, 8),
    to_signed(-28, 8),
    to_signed(-32, 8),
    to_signed(-30, 8),
    to_signed(-22, 8),
    to_signed(-10, 8),
    to_signed(4, 8),
    to_signed(17, 8),
    to_signed(25, 8),
    to_signed(30, 8),
    to_signed(33, 8),
    to_signed(33, 8),
    to_signed(30, 8),
    to_signed(26, 8),
    to_signed(20, 8),
    to_signed(13, 8),
    to_signed(7, 8),
    to_signed(2, 8),
    to_signed(-3, 8),
    to_signed(-8, 8),
    to_signed(-11, 8),
    to_signed(-8, 8),
    to_signed(2, 8),
    to_signed(18, 8),
    to_signed(36, 8),
    to_signed(52, 8),
    to_signed(62, 8),
    to_signed(65, 8),
    to_signed(61, 8),
    to_signed(53, 8),
    to_signed(40, 8),
    to_signed(25, 8),
    to_signed(12, 8),
    to_signed(1, 8),
    to_signed(-15, 8),
    to_signed(-37, 8),
    to_signed(-59, 8),
    to_signed(-69, 8),
    to_signed(-62, 8),
    to_signed(-41, 8),
    to_signed(-15, 8),
    to_signed(9, 8),
    to_signed(21, 8),
    to_signed(18, 8),
    to_signed(2, 8),
    to_signed(-25, 8),
    to_signed(-54, 8),
    to_signed(-76, 8),
    to_signed(-82, 8),
    to_signed(-71, 8),
    to_signed(-51, 8),
    to_signed(-25, 8),
    to_signed(6, 8),
    to_signed(37, 8),
    to_signed(61, 8),
    to_signed(74, 8),
    to_signed(77, 8),
    to_signed(72, 8),
    to_signed(59, 8),
    to_signed(42, 8),
    to_signed(27, 8),
    to_signed(16, 8),
    to_signed(8, 8),
    to_signed(3, 8),
    to_signed(-3, 8),
    to_signed(-10, 8),
    to_signed(-19, 8),
    to_signed(-23, 8),
    to_signed(-21, 8),
    to_signed(-17, 8),
    to_signed(-15, 8),
    to_signed(-12, 8),
    to_signed(-10, 8),
    to_signed(-11, 8),
    to_signed(-19, 8),
    to_signed(-29, 8),
    to_signed(-38, 8),
    to_signed(-42, 8),
    to_signed(-38, 8),
    to_signed(-24, 8),
    to_signed(-4, 8),
    to_signed(17, 8),
    to_signed(31, 8),
    to_signed(39, 8),
    to_signed(41, 8),
    to_signed(40, 8),
    to_signed(39, 8),
    to_signed(38, 8),
    to_signed(35, 8),
    to_signed(29, 8),
    to_signed(21, 8),
    to_signed(14, 8),
    to_signed(7, 8),
    to_signed(1, 8),
    to_signed(-4, 8),
    to_signed(-3, 8),
    to_signed(3, 8),
    to_signed(15, 8),
    to_signed(33, 8),
    to_signed(52, 8),
    to_signed(68, 8),
    to_signed(77, 8),
    to_signed(79, 8),
    to_signed(74, 8),
    to_signed(65, 8),
    to_signed(51, 8),
    to_signed(35, 8),
    to_signed(21, 8),
    to_signed(8, 8),
    to_signed(-8, 8),
    to_signed(-29, 8),
    to_signed(-52, 8),
    to_signed(-67, 8),
    to_signed(-65, 8),
    to_signed(-49, 8),
    to_signed(-27, 8),
    to_signed(-6, 8),
    to_signed(6, 8),
    to_signed(6, 8),
    to_signed(-6, 8),
    to_signed(-29, 8),
    to_signed(-55, 8),
    to_signed(-74, 8),
    to_signed(-78, 8),
    to_signed(-69, 8),
    to_signed(-50, 8),
    to_signed(-26, 8),
    to_signed(2, 8),
    to_signed(32, 8),
    to_signed(56, 8),
    to_signed(69, 8),
    to_signed(71, 8),
    to_signed(65, 8),
    to_signed(51, 8),
    to_signed(33, 8),
    to_signed(16, 8),
    to_signed(3, 8),
    to_signed(-5, 8),
    to_signed(-11, 8),
    to_signed(-15, 8),
    to_signed(-20, 8),
    to_signed(-25, 8),
    to_signed(-26, 8),
    to_signed(-20, 8),
    to_signed(-11, 8),
    to_signed(-5, 8),
    to_signed(-4, 8),
    to_signed(-5, 8),
    to_signed(-10, 8),
    to_signed(-18, 8),
    to_signed(-26, 8),
    to_signed(-31, 8),
    to_signed(-33, 8),
    to_signed(-29, 8),
    to_signed(-17, 8),
    to_signed(2, 8),
    to_signed(23, 8),
    to_signed(36, 8),
    to_signed(40, 8),
    to_signed(42, 8),
    to_signed(43, 8),
    to_signed(45, 8),
    to_signed(46, 8),
    to_signed(45, 8),
    to_signed(39, 8),
    to_signed(30, 8),
    to_signed(20, 8),
    to_signed(11, 8),
    to_signed(3, 8),
    to_signed(-2, 8),
    to_signed(-2, 8),
    to_signed(3, 8),
    to_signed(12, 8),
    to_signed(24, 8),
    to_signed(38, 8),
    to_signed(50, 8),
    to_signed(57, 8),
    to_signed(56, 8),
    to_signed(51, 8),
    to_signed(43, 8),
    to_signed(31, 8),
    to_signed(18, 8),
    to_signed(7, 8),
    to_signed(-4, 8),
    to_signed(-19, 8),
    to_signed(-40, 8),
    to_signed(-61, 8),
    to_signed(-72, 8),
    to_signed(-70, 8),
    to_signed(-55, 8),
    to_signed(-33, 8),
    to_signed(-13, 8),
    to_signed(-3, 8),
    to_signed(-4, 8),
    to_signed(-16, 8),
    to_signed(-38, 8),
    to_signed(-63, 8),
    to_signed(-83, 8),
    to_signed(-88, 8),
    to_signed(-81, 8),
    to_signed(-66, 8),
    to_signed(-46, 8),
    to_signed(-20, 8),
    to_signed(7, 8),
    to_signed(29, 8),
    to_signed(41, 8),
    to_signed(46, 8),
    to_signed(45, 8),
    to_signed(41, 8),
    to_signed(33, 8),
    to_signed(23, 8),
    to_signed(12, 8),
    to_signed(3, 8),
    to_signed(-6, 8),
    to_signed(-15, 8),
    to_signed(-25, 8),
    to_signed(-35, 8),
    to_signed(-39, 8),
    to_signed(-34, 8),
    to_signed(-24, 8),
    to_signed(-14, 8),
    to_signed(-8, 8),
    to_signed(-11, 8),
    to_signed(-19, 8),
    to_signed(-30, 8),
    to_signed(-40, 8),
    to_signed(-47, 8),
    to_signed(-49, 8),
    to_signed(-46, 8),
    to_signed(-34, 8),
    to_signed(-14, 8),
    to_signed(7, 8),
    to_signed(23, 8),
    to_signed(30, 8),
    to_signed(31, 8),
    to_signed(29, 8),
    to_signed(28, 8),
    to_signed(27, 8),
    to_signed(25, 8),
    to_signed(22, 8),
    to_signed(18, 8),
    to_signed(12, 8),
    to_signed(2, 8),
    to_signed(-10, 8),
    to_signed(-19, 8),
    to_signed(-21, 8),
    to_signed(-16, 8),
    to_signed(-4, 8),
    to_signed(11, 8),
    to_signed(27, 8),
    to_signed(43, 8),
    to_signed(53, 8),
    to_signed(57, 8),
    to_signed(56, 8),
    to_signed(49, 8),
    to_signed(39, 8),
    to_signed(25, 8),
    to_signed(10, 8),
    to_signed(-6, 8),
    to_signed(-27, 8),
    to_signed(-51, 8),
    to_signed(-74, 8),
    to_signed(-84, 8),
    to_signed(-78, 8),
    to_signed(-60, 8),
    to_signed(-37, 8),
    to_signed(-17, 8),
    to_signed(-7, 8),
    to_signed(-10, 8),
    to_signed(-25, 8),
    to_signed(-50, 8),
    to_signed(-75, 8),
    to_signed(-93, 8),
    to_signed(-97, 8),
    to_signed(-87, 8),
    to_signed(-69, 8),
    to_signed(-45, 8),
    to_signed(-16, 8),
    to_signed(15, 8),
    to_signed(38, 8),
    to_signed(50, 8),
    to_signed(51, 8),
    to_signed(46, 8),
    to_signed(37, 8),
    to_signed(25, 8),
    to_signed(12, 8),
    to_signed(-1, 8),
    to_signed(-12, 8),
    to_signed(-23, 8),
    to_signed(-32, 8),
    to_signed(-39, 8),
    to_signed(-43, 8),
    to_signed(-44, 8),
    to_signed(-38, 8),
    to_signed(-27, 8),
    to_signed(-16, 8),
    to_signed(-10, 8),
    to_signed(-12, 8),
    to_signed(-21, 8),
    to_signed(-32, 8),
    to_signed(-40, 8),
    to_signed(-40, 8),
    to_signed(-36, 8),
    to_signed(-27, 8),
    to_signed(-14, 8),
    to_signed(4, 8),
    to_signed(22, 8),
    to_signed(32, 8),
    to_signed(34, 8),
    to_signed(32, 8),
    to_signed(30, 8),
    to_signed(30, 8),
    to_signed(29, 8),
    to_signed(28, 8),
    to_signed(27, 8),
    to_signed(24, 8),
    to_signed(18, 8),
    to_signed(8, 8),
    to_signed(-5, 8),
    to_signed(-15, 8),
    to_signed(-17, 8),
    to_signed(-9, 8),
    to_signed(7, 8),
    to_signed(26, 8),
    to_signed(44, 8),
    to_signed(57, 8),
    to_signed(63, 8),
    to_signed(59, 8),
    to_signed(49, 8),
    to_signed(36, 8),
    to_signed(22, 8),
    to_signed(9, 8),
    to_signed(-1, 8),
    to_signed(-9, 8),
    to_signed(-21, 8),
    to_signed(-38, 8),
    to_signed(-56, 8),
    to_signed(-66, 8),
    to_signed(-63, 8),
    to_signed(-48, 8),
    to_signed(-29, 8),
    to_signed(-13, 8),
    to_signed(-2, 8),
    to_signed(-2, 8),
    to_signed(-13, 8),
    to_signed(-34, 8),
    to_signed(-57, 8),
    to_signed(-73, 8),
    to_signed(-76, 8),
    to_signed(-68, 8),
    to_signed(-52, 8),
    to_signed(-32, 8),
    to_signed(-8, 8),
    to_signed(16, 8),
    to_signed(35, 8),
    to_signed(44, 8),
    to_signed(44, 8),
    to_signed(39, 8),
    to_signed(32, 8),
    to_signed(25, 8),
    to_signed(18, 8),
    to_signed(13, 8),
    to_signed(7, 8),
    to_signed(-1, 8),
    to_signed(-9, 8),
    to_signed(-15, 8),
    to_signed(-19, 8),
    to_signed(-19, 8),
    to_signed(-15, 8),
    to_signed(-8, 8),
    to_signed(1, 8),
    to_signed(6, 8),
    to_signed(3, 8),
    to_signed(-6, 8),
    to_signed(-18, 8),
    to_signed(-28, 8),
    to_signed(-32, 8),
    to_signed(-30, 8),
    to_signed(-23, 8),
    to_signed(-13, 8),
    to_signed(3, 8),
    to_signed(20, 8),
    to_signed(32, 8),
    to_signed(37, 8),
    to_signed(37, 8),
    to_signed(37, 8),
    to_signed(38, 8),
    to_signed(38, 8),
    to_signed(36, 8),
    to_signed(34, 8),
    to_signed(33, 8),
    to_signed(31, 8),
    to_signed(26, 8),
    to_signed(19, 8),
    to_signed(11, 8),
    to_signed(7, 8),
    to_signed(11, 8),
    to_signed(22, 8),
    to_signed(37, 8),
    to_signed(51, 8),
    to_signed(62, 8),
    to_signed(68, 8),
    to_signed(65, 8),
    to_signed(58, 8),
    to_signed(49, 8),
    to_signed(41, 8),
    to_signed(33, 8),
    to_signed(24, 8),
    to_signed(14, 8),
    to_signed(-3, 8),
    to_signed(-26, 8),
    to_signed(-49, 8),
    to_signed(-60, 8),
    to_signed(-53, 8),
    to_signed(-33, 8),
    to_signed(-9, 8),
    to_signed(13, 8),
    to_signed(25, 8),
    to_signed(23, 8),
    to_signed(8, 8),
    to_signed(-18, 8),
    to_signed(-45, 8),
    to_signed(-65, 8),
    to_signed(-70, 8),
    to_signed(-59, 8),
    to_signed(-38, 8),
    to_signed(-14, 8),
    to_signed(11, 8),
    to_signed(35, 8),
    to_signed(53, 8),
    to_signed(62, 8),
    to_signed(65, 8),
    to_signed(61, 8),
    to_signed(53, 8),
    to_signed(41, 8),
    to_signed(30, 8),
    to_signed(21, 8),
    to_signed(13, 8),
    to_signed(5, 8),
    to_signed(-4, 8),
    to_signed(-13, 8),
    to_signed(-19, 8),
    to_signed(-20, 8),
    to_signed(-17, 8),
    to_signed(-12, 8),
    to_signed(-6, 8),
    to_signed(-2, 8),
    to_signed(-3, 8),
    to_signed(-10, 8),
    to_signed(-22, 8),
    to_signed(-31, 8),
    to_signed(-34, 8),
    to_signed(-29, 8),
    to_signed(-18, 8),
    to_signed(-3, 8),
    to_signed(15, 8),
    to_signed(32, 8),
    to_signed(43, 8),
    to_signed(46, 8),
    to_signed(43, 8),
    to_signed(41, 8),
    to_signed(41, 8),
    to_signed(44, 8),
    to_signed(47, 8),
    to_signed(48, 8),
    to_signed(46, 8),
    to_signed(39, 8),
    to_signed(26, 8),
    to_signed(10, 8),
    to_signed(-4, 8),
    to_signed(-9, 8),
    to_signed(-3, 8),
    to_signed(14, 8),
    to_signed(37, 8),
    to_signed(59, 8),
    to_signed(74, 8),
    to_signed(77, 8),
    to_signed(71, 8),
    to_signed(57, 8),
    to_signed(41, 8),
    to_signed(26, 8),
    to_signed(12, 8),
    to_signed(-1, 8),
    to_signed(-15, 8),
    to_signed(-33, 8),
    to_signed(-54, 8),
    to_signed(-71, 8),
    to_signed(-75, 8),
    to_signed(-62, 8),
    to_signed(-38, 8),
    to_signed(-13, 8),
    to_signed(3, 8),
    to_signed(8, 8),
    to_signed(0, 8),
    to_signed(-19, 8),
    to_signed(-44, 8),
    to_signed(-67, 8),
    to_signed(-82, 8),
    to_signed(-83, 8),
    to_signed(-70, 8),
    to_signed(-48, 8),
    to_signed(-21, 8),
    to_signed(5, 8),
    to_signed(26, 8),
    to_signed(40, 8),
    to_signed(46, 8),
    to_signed(44, 8),
    to_signed(39, 8),
    to_signed(32, 8),
    to_signed(23, 8),
    to_signed(12, 8),
    to_signed(4, 8),
    to_signed(-3, 8),
    to_signed(-11, 8),
    to_signed(-21, 8),
    to_signed(-32, 8),
    to_signed(-40, 8),
    to_signed(-39, 8),
    to_signed(-30, 8),
    to_signed(-14, 8),
    to_signed(1, 8),
    to_signed(11, 8),
    to_signed(11, 8),
    to_signed(3, 8),
    to_signed(-11, 8),
    to_signed(-25, 8),
    to_signed(-33, 8),
    to_signed(-32, 8),
    to_signed(-23, 8),
    to_signed(-9, 8),
    to_signed(8, 8),
    to_signed(22, 8),
    to_signed(31, 8),
    to_signed(33, 8),
    to_signed(34, 8),
    to_signed(34, 8),
    to_signed(34, 8),
    to_signed(34, 8),
    to_signed(34, 8),
    to_signed(32, 8),
    to_signed(26, 8),
    to_signed(15, 8),
    to_signed(1, 8),
    to_signed(-13, 8),
    to_signed(-21, 8),
    to_signed(-21, 8),
    to_signed(-11, 8),
    to_signed(6, 8),
    to_signed(26, 8),
    to_signed(45, 8),
    to_signed(57, 8),
    to_signed(58, 8),
    to_signed(49, 8),
    to_signed(33, 8),
    to_signed(17, 8),
    to_signed(4, 8),
    to_signed(-7, 8),
    to_signed(-18, 8),
    to_signed(-29, 8),
    to_signed(-44, 8),
    to_signed(-61, 8),
    to_signed(-76, 8),
    to_signed(-79, 8),
    to_signed(-68, 8),
    to_signed(-45, 8),
    to_signed(-21, 8),
    to_signed(-4, 8),
    to_signed(1, 8),
    to_signed(-4, 8),
    to_signed(-18, 8),
    to_signed(-38, 8),
    to_signed(-59, 8),
    to_signed(-76, 8),
    to_signed(-83, 8),
    to_signed(-79, 8),
    to_signed(-65, 8),
    to_signed(-42, 8),
    to_signed(-14, 8),
    to_signed(12, 8),
    to_signed(32, 8),
    to_signed(44, 8),
    to_signed(48, 8),
    to_signed(47, 8),
    to_signed(44, 8),
    to_signed(37, 8),
    to_signed(27, 8),
    to_signed(15, 8),
    to_signed(3, 8),
    to_signed(-8, 8),
    to_signed(-20, 8),
    to_signed(-32, 8),
    to_signed(-41, 8),
    to_signed(-41, 8),
    to_signed(-31, 8),
    to_signed(-13, 8),
    to_signed(4, 8),
    to_signed(13, 8),
    to_signed(9, 8),
    to_signed(-6, 8),
    to_signed(-26, 8),
    to_signed(-45, 8),
    to_signed(-56, 8),
    to_signed(-57, 8),
    to_signed(-47, 8),
    to_signed(-31, 8),
    to_signed(-13, 8),
    to_signed(2, 8),
    to_signed(11, 8),
    to_signed(16, 8),
    to_signed(20, 8),
    to_signed(24, 8),
    to_signed(27, 8),
    to_signed(27, 8),
    to_signed(26, 8),
    to_signed(23, 8),
    to_signed(18, 8),
    to_signed(8, 8),
    to_signed(-7, 8),
    to_signed(-22, 8),
    to_signed(-31, 8),
    to_signed(-31, 8),
    to_signed(-21, 8),
    to_signed(-4, 8),
    to_signed(16, 8),
    to_signed(36, 8),
    to_signed(52, 8),
    to_signed(60, 8),
    to_signed(56, 8),
    to_signed(43, 8),
    to_signed(27, 8),
    to_signed(12, 8),
    to_signed(-1, 8),
    to_signed(-13, 8),
    to_signed(-28, 8),
    to_signed(-45, 8),
    to_signed(-63, 8),
    to_signed(-77, 8),
    to_signed(-81, 8),
    to_signed(-71, 8),
    to_signed(-51, 8),
    to_signed(-29, 8),
    to_signed(-13, 8),
    to_signed(-8, 8),
    to_signed(-15, 8),
    to_signed(-31, 8),
    to_signed(-51, 8),
    to_signed(-68, 8),
    to_signed(-80, 8),
    to_signed(-83, 8),
    to_signed(-78, 8),
    to_signed(-66, 8),
    to_signed(-45, 8),
    to_signed(-20, 8),
    to_signed(7, 8),
    to_signed(30, 8),
    to_signed(45, 8),
    to_signed(53, 8),
    to_signed(54, 8),
    to_signed(51, 8),
    to_signed(44, 8),
    to_signed(34, 8),
    to_signed(22, 8),
    to_signed(8, 8),
    to_signed(-6, 8),
    to_signed(-19, 8),
    to_signed(-32, 8),
    to_signed(-41, 8),
    to_signed(-44, 8),
    to_signed(-36, 8),
    to_signed(-21, 8),
    to_signed(-5, 8),
    to_signed(6, 8),
    to_signed(6, 8),
    to_signed(-4, 8),
    to_signed(-21, 8),
    to_signed(-35, 8),
    to_signed(-43, 8),
    to_signed(-42, 8),
    to_signed(-34, 8),
    to_signed(-19, 8),
    to_signed(-3, 8),
    to_signed(9, 8),
    to_signed(15, 8),
    to_signed(18, 8),
    to_signed(21, 8),
    to_signed(27, 8),
    to_signed(36, 8),
    to_signed(42, 8),
    to_signed(44, 8),
    to_signed(43, 8),
    to_signed(38, 8),
    to_signed(28, 8),
    to_signed(12, 8),
    to_signed(-6, 8),
    to_signed(-18, 8),
    to_signed(-19, 8),
    to_signed(-10, 8),
    to_signed(8, 8),
    to_signed(28, 8),
    to_signed(47, 8),
    to_signed(61, 8),
    to_signed(69, 8),
    to_signed(69, 8),
    to_signed(59, 8),
    to_signed(44, 8),
    to_signed(29, 8),
    to_signed(16, 8),
    to_signed(3, 8),
    to_signed(-16, 8),
    to_signed(-41, 8),
    to_signed(-67, 8),
    to_signed(-86, 8),
    to_signed(-89, 8),
    to_signed(-76, 8),
    to_signed(-50, 8),
    to_signed(-19, 8),
    to_signed(6, 8),
    to_signed(19, 8),
    to_signed(17, 8),
    to_signed(0, 8),
    to_signed(-25, 8),
    to_signed(-50, 8),
    to_signed(-67, 8),
    to_signed(-72, 8),
    to_signed(-69, 8),
    to_signed(-57, 8),
    to_signed(-37, 8),
    to_signed(-11, 8),
    to_signed(15, 8),
    to_signed(38, 8),
    to_signed(55, 8),
    to_signed(66, 8),
    to_signed(70, 8),
    to_signed(67, 8),
    to_signed(59, 8),
    to_signed(48, 8),
    to_signed(36, 8),
    to_signed(24, 8),
    to_signed(9, 8),
    to_signed(-7, 8),
    to_signed(-22, 8),
    to_signed(-32, 8),
    to_signed(-34, 8),
    to_signed(-27, 8),
    to_signed(-13, 8),
    to_signed(1, 8),
    to_signed(10, 8),
    to_signed(9, 8),
    to_signed(-2, 8),
    to_signed(-18, 8),
    to_signed(-34, 8),
    to_signed(-44, 8),
    to_signed(-45, 8),
    to_signed(-39, 8),
    to_signed(-29, 8),
    to_signed(-15, 8),
    to_signed(0, 8),
    to_signed(12, 8),
    to_signed(20, 8),
    to_signed(26, 8),
    to_signed(33, 8),
    to_signed(42, 8),
    to_signed(51, 8),
    to_signed(56, 8),
    to_signed(54, 8),
    to_signed(47, 8),
    to_signed(34, 8),
    to_signed(17, 8),
    to_signed(-4, 8),
    to_signed(-20, 8),
    to_signed(-25, 8),
    to_signed(-16, 8),
    to_signed(5, 8),
    to_signed(33, 8),
    to_signed(59, 8),
    to_signed(76, 8),
    to_signed(82, 8),
    to_signed(79, 8),
    to_signed(68, 8),
    to_signed(50, 8),
    to_signed(33, 8),
    to_signed(20, 8),
    to_signed(12, 8),
    to_signed(0, 8),
    to_signed(-20, 8),
    to_signed(-46, 8),
    to_signed(-67, 8),
    to_signed(-72, 8),
    to_signed(-60, 8),
    to_signed(-35, 8),
    to_signed(-7, 8),
    to_signed(16, 8),
    to_signed(26, 8),
    to_signed(21, 8),
    to_signed(0, 8),
    to_signed(-30, 8),
    to_signed(-58, 8),
    to_signed(-76, 8),
    to_signed(-80, 8),
    to_signed(-70, 8),
    to_signed(-51, 8),
    to_signed(-29, 8),
    to_signed(-5, 8),
    to_signed(18, 8),
    to_signed(34, 8),
    to_signed(44, 8),
    to_signed(49, 8),
    to_signed(51, 8),
    to_signed(49, 8),
    to_signed(40, 8),
    to_signed(28, 8),
    to_signed(16, 8),
    to_signed(6, 8),
    to_signed(-6, 8),
    to_signed(-21, 8),
    to_signed(-37, 8),
    to_signed(-50, 8),
    to_signed(-53, 8),
    to_signed(-46, 8),
    to_signed(-34, 8),
    to_signed(-20, 8),
    to_signed(-10, 8),
    to_signed(-8, 8),
    to_signed(-14, 8),
    to_signed(-25, 8),
    to_signed(-34, 8),
    to_signed(-37, 8),
    to_signed(-34, 8),
    to_signed(-26, 8),
    to_signed(-16, 8),
    to_signed(-4, 8),
    to_signed(9, 8),
    to_signed(23, 8),
    to_signed(35, 8),
    to_signed(41, 8),
    to_signed(42, 8),
    to_signed(45, 8),
    to_signed(50, 8),
    to_signed(56, 8),
    to_signed(56, 8),
    to_signed(50, 8),
    to_signed(38, 8),
    to_signed(22, 8),
    to_signed(4, 8),
    to_signed(-11, 8),
    to_signed(-16, 8),
    to_signed(-8, 8),
    to_signed(14, 8),
    to_signed(42, 8),
    to_signed(69, 8),
    to_signed(86, 8),
    to_signed(90, 8),
    to_signed(83, 8),
    to_signed(67, 8),
    to_signed(47, 8),
    to_signed(28, 8),
    to_signed(16, 8),
    to_signed(10, 8),
    to_signed(3, 8),
    to_signed(-13, 8),
    to_signed(-39, 8),
    to_signed(-67, 8),
    to_signed(-83, 8),
    to_signed(-79, 8),
    to_signed(-57, 8),
    to_signed(-29, 8),
    to_signed(-3, 8),
    to_signed(14, 8),
    to_signed(17, 8),
    to_signed(4, 8),
    to_signed(-22, 8),
    to_signed(-50, 8),
    to_signed(-73, 8),
    to_signed(-84, 8),
    to_signed(-80, 8),
    to_signed(-63, 8),
    to_signed(-38, 8),
    to_signed(-9, 8),
    to_signed(19, 8),
    to_signed(43, 8),
    to_signed(56, 8),
    to_signed(59, 8),
    to_signed(57, 8),
    to_signed(50, 8),
    to_signed(39, 8),
    to_signed(25, 8),
    to_signed(13, 8),
    to_signed(6, 8),
    to_signed(3, 8),
    to_signed(-1, 8),
    to_signed(-8, 8),
    to_signed(-17, 8),
    to_signed(-23, 8),
    to_signed(-20, 8),
    to_signed(-9, 8),
    to_signed(5, 8),
    to_signed(17, 8),
    to_signed(20, 8),
    to_signed(13, 8),
    to_signed(-3, 8),
    to_signed(-20, 8),
    to_signed(-29, 8),
    to_signed(-28, 8),
    to_signed(-18, 8),
    to_signed(-3, 8),
    to_signed(12, 8),
    to_signed(24, 8),
    to_signed(34, 8),
    to_signed(43, 8),
    to_signed(48, 8),
    to_signed(46, 8),
    to_signed(41, 8),
    to_signed(39, 8),
    to_signed(42, 8),
    to_signed(43, 8),
    to_signed(40, 8),
    to_signed(29, 8),
    to_signed(15, 8),
    to_signed(-1, 8),
    to_signed(-12, 8),
    to_signed(-18, 8),
    to_signed(-16, 8),
    to_signed(-4, 8),
    to_signed(17, 8),
    to_signed(38, 8),
    to_signed(55, 8),
    to_signed(63, 8),
    to_signed(60, 8),
    to_signed(49, 8),
    to_signed(31, 8),
    to_signed(14, 8),
    to_signed(2, 8),
    to_signed(-2, 8),
    to_signed(-1, 8),
    to_signed(-2, 8),
    to_signed(-13, 8),
    to_signed(-35, 8),
    to_signed(-56, 8),
    to_signed(-66, 8),
    to_signed(-61, 8),
    to_signed(-45, 8),
    to_signed(-24, 8),
    to_signed(-4, 8),
    to_signed(8, 8),
    to_signed(6, 8),
    to_signed(-9, 8),
    to_signed(-33, 8),
    to_signed(-57, 8),
    to_signed(-74, 8),
    to_signed(-79, 8),
    to_signed(-70, 8),
    to_signed(-50, 8),
    to_signed(-22, 8),
    to_signed(9, 8),
    to_signed(34, 8),
    to_signed(51, 8),
    to_signed(56, 8),
    to_signed(52, 8),
    to_signed(42, 8),
    to_signed(30, 8),
    to_signed(18, 8),
    to_signed(7, 8),
    to_signed(-2, 8),
    to_signed(-7, 8),
    to_signed(-9, 8),
    to_signed(-13, 8),
    to_signed(-22, 8),
    to_signed(-31, 8),
    to_signed(-37, 8),
    to_signed(-36, 8),
    to_signed(-29, 8),
    to_signed(-21, 8),
    to_signed(-15, 8),
    to_signed(-17, 8),
    to_signed(-26, 8),
    to_signed(-37, 8),
    to_signed(-45, 8),
    to_signed(-44, 8),
    to_signed(-36, 8),
    to_signed(-23, 8),
    to_signed(-8, 8),
    to_signed(5, 8),
    to_signed(14, 8),
    to_signed(21, 8),
    to_signed(26, 8),
    to_signed(28, 8),
    to_signed(25, 8),
    to_signed(20, 8),
    to_signed(19, 8),
    to_signed(20, 8),
    to_signed(21, 8),
    to_signed(16, 8),
    to_signed(6, 8),
    to_signed(-5, 8),
    to_signed(-15, 8),
    to_signed(-23, 8),
    to_signed(-28, 8),
    to_signed(-25, 8),
    to_signed(-14, 8),
    to_signed(5, 8),
    to_signed(27, 8),
    to_signed(45, 8),
    to_signed(56, 8),
    to_signed(56, 8),
    to_signed(49, 8),
    to_signed(37, 8),
    to_signed(25, 8),
    to_signed(17, 8),
    to_signed(14, 8),
    to_signed(13, 8),
    to_signed(7, 8),
    to_signed(-8, 8),
    to_signed(-32, 8),
    to_signed(-55, 8),
    to_signed(-68, 8),
    to_signed(-65, 8),
    to_signed(-50, 8),
    to_signed(-28, 8),
    to_signed(-9, 8),
    to_signed(0, 8),
    to_signed(-5, 8),
    to_signed(-21, 8),
    to_signed(-45, 8),
    to_signed(-66, 8),
    to_signed(-80, 8),
    to_signed(-82, 8),
    to_signed(-71, 8),
    to_signed(-49, 8),
    to_signed(-22, 8),
    to_signed(5, 8),
    to_signed(27, 8),
    to_signed(43, 8),
    to_signed(50, 8),
    to_signed(48, 8),
    to_signed(41, 8),
    to_signed(29, 8),
    to_signed(15, 8),
    to_signed(-1, 8),
    to_signed(-12, 8),
    to_signed(-14, 8),
    to_signed(-10, 8),
    to_signed(-6, 8),
    to_signed(-5, 8),
    to_signed(-8, 8),
    to_signed(-12, 8),
    to_signed(-14, 8),
    to_signed(-11, 8),
    to_signed(-7, 8),
    to_signed(-5, 8),
    to_signed(-6, 8),
    to_signed(-10, 8),
    to_signed(-15, 8),
    to_signed(-21, 8),
    to_signed(-22, 8),
    to_signed(-18, 8),
    to_signed(-11, 8),
    to_signed(0, 8),
    to_signed(13, 8),
    to_signed(25, 8),
    to_signed(34, 8),
    to_signed(40, 8),
    to_signed(41, 8),
    to_signed(38, 8),
    to_signed(34, 8),
    to_signed(34, 8),
    to_signed(37, 8),
    to_signed(37, 8),
    to_signed(33, 8),
    to_signed(29, 8),
    to_signed(25, 8),
    to_signed(21, 8),
    to_signed(15, 8),
    to_signed(11, 8),
    to_signed(12, 8),
    to_signed(18, 8),
    to_signed(29, 8),
    to_signed(44, 8),
    to_signed(57, 8),
    to_signed(62, 8),
    to_signed(61, 8),
    to_signed(56, 8),
    to_signed(48, 8),
    to_signed(38, 8),
    to_signed(31, 8),
    to_signed(25, 8),
    to_signed(18, 8),
    to_signed(7, 8),
    to_signed(-11, 8),
    to_signed(-36, 8),
    to_signed(-61, 8),
    to_signed(-75, 8),
    to_signed(-69, 8),
    to_signed(-48, 8),
    to_signed(-24, 8),
    to_signed(-3, 8),
    to_signed(7, 8),
    to_signed(3, 8),
    to_signed(-14, 8),
    to_signed(-36, 8),
    to_signed(-57, 8),
    to_signed(-71, 8),
    to_signed(-73, 8),
    to_signed(-61, 8),
    to_signed(-40, 8),
    to_signed(-17, 8),
    to_signed(5, 8),
    to_signed(27, 8),
    to_signed(42, 8),
    to_signed(48, 8),
    to_signed(47, 8),
    to_signed(42, 8),
    to_signed(31, 8),
    to_signed(18, 8),
    to_signed(5, 8),
    to_signed(-3, 8),
    to_signed(-5, 8),
    to_signed(-3, 8),
    to_signed(-2, 8),
    to_signed(-5, 8),
    to_signed(-13, 8),
    to_signed(-21, 8),
    to_signed(-21, 8),
    to_signed(-17, 8),
    to_signed(-12, 8),
    to_signed(-10, 8),
    to_signed(-12, 8),
    to_signed(-19, 8),
    to_signed(-27, 8),
    to_signed(-31, 8),
    to_signed(-30, 8),
    to_signed(-26, 8),
    to_signed(-18, 8),
    to_signed(-6, 8),
    to_signed(9, 8),
    to_signed(21, 8),
    to_signed(29, 8),
    to_signed(33, 8),
    to_signed(33, 8),
    to_signed(29, 8),
    to_signed(25, 8),
    to_signed(24, 8),
    to_signed(24, 8),
    to_signed(21, 8),
    to_signed(17, 8),
    to_signed(15, 8),
    to_signed(13, 8),
    to_signed(8, 8),
    to_signed(1, 8),
    to_signed(-4, 8),
    to_signed(-5, 8),
    to_signed(-1, 8),
    to_signed(12, 8),
    to_signed(28, 8),
    to_signed(40, 8),
    to_signed(48, 8),
    to_signed(50, 8),
    to_signed(47, 8),
    to_signed(39, 8),
    to_signed(29, 8),
    to_signed(21, 8),
    to_signed(16, 8),
    to_signed(8, 8),
    to_signed(-4, 8),
    to_signed(-25, 8),
    to_signed(-53, 8),
    to_signed(-79, 8),
    to_signed(-89, 8),
    to_signed(-81, 8),
    to_signed(-62, 8),
    to_signed(-38, 8),
    to_signed(-18, 8),
    to_signed(-8, 8),
    to_signed(-13, 8),
    to_signed(-29, 8),
    to_signed(-50, 8),
    to_signed(-69, 8),
    to_signed(-81, 8),
    to_signed(-80, 8),
    to_signed(-65, 8),
    to_signed(-44, 8),
    to_signed(-21, 8),
    to_signed(3, 8),
    to_signed(24, 8),
    to_signed(38, 8),
    to_signed(43, 8),
    to_signed(43, 8),
    to_signed(38, 8),
    to_signed(29, 8),
    to_signed(16, 8),
    to_signed(5, 8),
    to_signed(-4, 8),
    to_signed(-10, 8),
    to_signed(-11, 8),
    to_signed(-11, 8),
    to_signed(-16, 8),
    to_signed(-23, 8),
    to_signed(-27, 8),
    to_signed(-24, 8),
    to_signed(-16, 8),
    to_signed(-8, 8),
    to_signed(-4, 8),
    to_signed(-6, 8),
    to_signed(-14, 8),
    to_signed(-23, 8),
    to_signed(-29, 8),
    to_signed(-32, 8),
    to_signed(-31, 8),
    to_signed(-24, 8),
    to_signed(-9, 8),
    to_signed(10, 8),
    to_signed(25, 8),
    to_signed(35, 8),
    to_signed(38, 8),
    to_signed(33, 8),
    to_signed(25, 8),
    to_signed(18, 8),
    to_signed(14, 8),
    to_signed(11, 8),
    to_signed(10, 8),
    to_signed(11, 8),
    to_signed(12, 8),
    to_signed(11, 8),
    to_signed(9, 8),
    to_signed(6, 8),
    to_signed(4, 8),
    to_signed(4, 8),
    to_signed(6, 8),
    to_signed(12, 8),
    to_signed(20, 8),
    to_signed(30, 8),
    to_signed(38, 8),
    to_signed(43, 8),
    to_signed(43, 8),
    to_signed(39, 8),
    to_signed(32, 8),
    to_signed(24, 8),
    to_signed(16, 8),
    to_signed(5, 8),
    to_signed(-10, 8),
    to_signed(-32, 8),
    to_signed(-58, 8),
    to_signed(-78, 8),
    to_signed(-84, 8),
    to_signed(-72, 8),
    to_signed(-50, 8),
    to_signed(-23, 8),
    to_signed(-3, 8),
    to_signed(4, 8),
    to_signed(-4, 8),
    to_signed(-24, 8),
    to_signed(-48, 8),
    to_signed(-67, 8),
    to_signed(-75, 8),
    to_signed(-68, 8),
    to_signed(-49, 8),
    to_signed(-23, 8),
    to_signed(4, 8),
    to_signed(28, 8),
    to_signed(47, 8),
    to_signed(58, 8),
    to_signed(61, 8),
    to_signed(59, 8),
    to_signed(54, 8),
    to_signed(46, 8),
    to_signed(35, 8),
    to_signed(22, 8),
    to_signed(12, 8),
    to_signed(9, 8),
    to_signed(10, 8),
    to_signed(10, 8),
    to_signed(4, 8),
    to_signed(-4, 8),
    to_signed(-10, 8),
    to_signed(-10, 8),
    to_signed(-6, 8),
    to_signed(-2, 8),
    to_signed(-4, 8),
    to_signed(-11, 8),
    to_signed(-21, 8),
    to_signed(-28, 8),
    to_signed(-31, 8),
    to_signed(-28, 8),
    to_signed(-21, 8),
    to_signed(-8, 8),
    to_signed(8, 8),
    to_signed(24, 8),
    to_signed(34, 8),
    to_signed(38, 8),
    to_signed(37, 8),
    to_signed(34, 8),
    to_signed(30, 8),
    to_signed(25, 8),
    to_signed(22, 8),
    to_signed(19, 8),
    to_signed(18, 8),
    to_signed(18, 8),
    to_signed(17, 8),
    to_signed(15, 8),
    to_signed(10, 8),
    to_signed(4, 8),
    to_signed(-3, 8),
    to_signed(-8, 8),
    to_signed(-10, 8),
    to_signed(-6, 8),
    to_signed(5, 8),
    to_signed(21, 8),
    to_signed(36, 8),
    to_signed(42, 8),
    to_signed(41, 8),
    to_signed(35, 8),
    to_signed(28, 8),
    to_signed(21, 8),
    to_signed(17, 8),
    to_signed(14, 8),
    to_signed(7, 8),
    to_signed(-8, 8),
    to_signed(-29, 8),
    to_signed(-50, 8),
    to_signed(-62, 8),
    to_signed(-58, 8),
    to_signed(-40, 8),
    to_signed(-21, 8),
    to_signed(-7, 8),
    to_signed(-4, 8),
    to_signed(-12, 8),
    to_signed(-28, 8),
    to_signed(-45, 8),
    to_signed(-57, 8),
    to_signed(-61, 8),
    to_signed(-55, 8),
    to_signed(-41, 8),
    to_signed(-21, 8),
    to_signed(-1, 8),
    to_signed(15, 8),
    to_signed(29, 8),
    to_signed(39, 8),
    to_signed(44, 8),
    to_signed(45, 8),
    to_signed(46, 8),
    to_signed(43, 8),
    to_signed(35, 8),
    to_signed(22, 8),
    to_signed(10, 8),
    to_signed(2, 8),
    to_signed(-4, 8),
    to_signed(-9, 8),
    to_signed(-17, 8),
    to_signed(-26, 8),
    to_signed(-31, 8),
    to_signed(-28, 8),
    to_signed(-20, 8),
    to_signed(-16, 8),
    to_signed(-18, 8),
    to_signed(-25, 8),
    to_signed(-35, 8),
    to_signed(-45, 8),
    to_signed(-49, 8),
    to_signed(-46, 8),
    to_signed(-37, 8),
    to_signed(-24, 8),
    to_signed(-7, 8),
    to_signed(9, 8),
    to_signed(20, 8),
    to_signed(25, 8),
    to_signed(27, 8),
    to_signed(24, 8),
    to_signed(17, 8),
    to_signed(10, 8),
    to_signed(7, 8),
    to_signed(8, 8),
    to_signed(13, 8),
    to_signed(20, 8),
    to_signed(25, 8),
    to_signed(26, 8),
    to_signed(23, 8),
    to_signed(16, 8),
    to_signed(9, 8),
    to_signed(4, 8),
    to_signed(3, 8),
    to_signed(9, 8),
    to_signed(19, 8),
    to_signed(33, 8),
    to_signed(45, 8),
    to_signed(53, 8),
    to_signed(53, 8),
    to_signed(49, 8),
    to_signed(42, 8),
    to_signed(36, 8),
    to_signed(30, 8),
    to_signed(24, 8),
    to_signed(17, 8),
    to_signed(3, 8),
    to_signed(-18, 8),
    to_signed(-41, 8),
    to_signed(-56, 8),
    to_signed(-55, 8),
    to_signed(-42, 8),
    to_signed(-23, 8),
    to_signed(-7, 8),
    to_signed(0, 8),
    to_signed(-2, 8),
    to_signed(-12, 8),
    to_signed(-24, 8),
    to_signed(-38, 8),
    to_signed(-48, 8),
    to_signed(-51, 8),
    to_signed(-45, 8),
    to_signed(-32, 8),
    to_signed(-17, 8),
    to_signed(0, 8),
    to_signed(16, 8),
    to_signed(28, 8),
    to_signed(34, 8),
    to_signed(38, 8),
    to_signed(40, 8),
    to_signed(40, 8),
    to_signed(35, 8),
    to_signed(24, 8),
    to_signed(11, 8),
    to_signed(0, 8),
    to_signed(-6, 8),
    to_signed(-9, 8),
    to_signed(-15, 8),
    to_signed(-24, 8),
    to_signed(-30, 8),
    to_signed(-28, 8),
    to_signed(-20, 8),
    to_signed(-14, 8),
    to_signed(-12, 8),
    to_signed(-15, 8),
    to_signed(-22, 8),
    to_signed(-30, 8),
    to_signed(-36, 8),
    to_signed(-35, 8),
    to_signed(-29, 8),
    to_signed(-17, 8),
    to_signed(-1, 8),
    to_signed(14, 8),
    to_signed(25, 8),
    to_signed(32, 8),
    to_signed(38, 8),
    to_signed(39, 8),
    to_signed(35, 8),
    to_signed(29, 8),
    to_signed(26, 8),
    to_signed(28, 8),
    to_signed(33, 8),
    to_signed(38, 8),
    to_signed(41, 8),
    to_signed(40, 8),
    to_signed(34, 8),
    to_signed(25, 8),
    to_signed(12, 8),
    to_signed(1, 8),
    to_signed(-4, 8),
    to_signed(-1, 8),
    to_signed(8, 8),
    to_signed(20, 8),
    to_signed(34, 8),
    to_signed(43, 8),
    to_signed(42, 8),
    to_signed(34, 8),
    to_signed(22, 8),
    to_signed(11, 8),
    to_signed(4, 8),
    to_signed(2, 8),
    to_signed(1, 8),
    to_signed(-5, 8),
    to_signed(-23, 8),
    to_signed(-48, 8),
    to_signed(-70, 8),
    to_signed(-80, 8),
    to_signed(-75, 8),
    to_signed(-56, 8),
    to_signed(-34, 8),
    to_signed(-20, 8),
    to_signed(-17, 8),
    to_signed(-20, 8),
    to_signed(-29, 8),
    to_signed(-42, 8),
    to_signed(-55, 8),
    to_signed(-62, 8),
    to_signed(-62, 8),
    to_signed(-52, 8),
    to_signed(-35, 8),
    to_signed(-14, 8),
    to_signed(8, 8),
    to_signed(27, 8),
    to_signed(42, 8),
    to_signed(51, 8),
    to_signed(55, 8),
    to_signed(56, 8),
    to_signed(51, 8),
    to_signed(39, 8),
    to_signed(22, 8),
    to_signed(7, 8),
    to_signed(-2, 8),
    to_signed(-7, 8),
    to_signed(-13, 8),
    to_signed(-22, 8),
    to_signed(-31, 8),
    to_signed(-35, 8),
    to_signed(-30, 8),
    to_signed(-23, 8),
    to_signed(-20, 8),
    to_signed(-23, 8),
    to_signed(-29, 8),
    to_signed(-36, 8),
    to_signed(-42, 8),
    to_signed(-45, 8),
    to_signed(-41, 8),
    to_signed(-30, 8),
    to_signed(-17, 8),
    to_signed(-4, 8),
    to_signed(7, 8),
    to_signed(16, 8),
    to_signed(23, 8),
    to_signed(24, 8),
    to_signed(19, 8),
    to_signed(9, 8),
    to_signed(1, 8),
    to_signed(0, 8),
    to_signed(5, 8),
    to_signed(12, 8),
    to_signed(16, 8),
    to_signed(18, 8),
    to_signed(16, 8),
    to_signed(9, 8),
    to_signed(-4, 8),
    to_signed(-17, 8),
    to_signed(-22, 8),
    to_signed(-18, 8),
    to_signed(-7, 8),
    to_signed(9, 8),
    to_signed(27, 8),
    to_signed(41, 8),
    to_signed(47, 8),
    to_signed(45, 8),
    to_signed(38, 8),
    to_signed(28, 8),
    to_signed(20, 8),
    to_signed(18, 8),
    to_signed(17, 8),
    to_signed(11, 8),
    to_signed(-6, 8),
    to_signed(-30, 8),
    to_signed(-54, 8),
    to_signed(-68, 8),
    to_signed(-66, 8),
    to_signed(-48, 8),
    to_signed(-23, 8),
    to_signed(-3, 8),
    to_signed(9, 8),
    to_signed(12, 8),
    to_signed(8, 8),
    to_signed(-5, 8),
    to_signed(-22, 8),
    to_signed(-39, 8),
    to_signed(-50, 8),
    to_signed(-48, 8),
    to_signed(-34, 8),
    to_signed(-11, 8),
    to_signed(15, 8),
    to_signed(41, 8),
    to_signed(60, 8),
    to_signed(69, 8),
    to_signed(69, 8),
    to_signed(66, 8),
    to_signed(59, 8),
    to_signed(46, 8),
    to_signed(28, 8),
    to_signed(12, 8),
    to_signed(1, 8),
    to_signed(-6, 8),
    to_signed(-12, 8),
    to_signed(-20, 8),
    to_signed(-30, 8),
    to_signed(-36, 8),
    to_signed(-33, 8),
    to_signed(-25, 8),
    to_signed(-19, 8),
    to_signed(-20, 8),
    to_signed(-26, 8),
    to_signed(-36, 8),
    to_signed(-49, 8),
    to_signed(-57, 8),
    to_signed(-57, 8),
    to_signed(-49, 8),
    to_signed(-36, 8),
    to_signed(-20, 8),
    to_signed(-3, 8),
    to_signed(11, 8),
    to_signed(22, 8),
    to_signed(28, 8),
    to_signed(27, 8),
    to_signed(20, 8),
    to_signed(14, 8),
    to_signed(15, 8),
    to_signed(21, 8),
    to_signed(27, 8),
    to_signed(30, 8),
    to_signed(31, 8),
    to_signed(28, 8),
    to_signed(19, 8),
    to_signed(7, 8),
    to_signed(-4, 8),
    to_signed(-9, 8),
    to_signed(-7, 8),
    to_signed(2, 8),
    to_signed(16, 8),
    to_signed(31, 8),
    to_signed(46, 8),
    to_signed(55, 8),
    to_signed(58, 8),
    to_signed(52, 8),
    to_signed(41, 8),
    to_signed(32, 8),
    to_signed(27, 8),
    to_signed(25, 8),
    to_signed(20, 8),
    to_signed(6, 8),
    to_signed(-17, 8),
    to_signed(-41, 8),
    to_signed(-59, 8),
    to_signed(-63, 8),
    to_signed(-51, 8),
    to_signed(-29, 8),
    to_signed(-7, 8),
    to_signed(8, 8),
    to_signed(10, 8),
    to_signed(-1, 8),
    to_signed(-21, 8),
    to_signed(-46, 8),
    to_signed(-67, 8),
    to_signed(-79, 8),
    to_signed(-76, 8),
    to_signed(-59, 8),
    to_signed(-32, 8),
    to_signed(0, 8),
    to_signed(29, 8),
    to_signed(51, 8),
    to_signed(60, 8),
    to_signed(62, 8),
    to_signed(60, 8),
    to_signed(55, 8),
    to_signed(45, 8),
    to_signed(30, 8),
    to_signed(15, 8),
    to_signed(5, 8),
    to_signed(-1, 8),
    to_signed(-5, 8),
    to_signed(-12, 8),
    to_signed(-23, 8),
    to_signed(-34, 8),
    to_signed(-38, 8),
    to_signed(-33, 8),
    to_signed(-25, 8),
    to_signed(-23, 8),
    to_signed(-27, 8),
    to_signed(-35, 8),
    to_signed(-45, 8),
    to_signed(-53, 8),
    to_signed(-55, 8),
    to_signed(-48, 8),
    to_signed(-33, 8),
    to_signed(-13, 8),
    to_signed(6, 8),
    to_signed(21, 8),
    to_signed(31, 8),
    to_signed(35, 8),
    to_signed(33, 8),
    to_signed(27, 8),
    to_signed(19, 8),
    to_signed(17, 8),
    to_signed(21, 8),
    to_signed(26, 8),
    to_signed(29, 8),
    to_signed(28, 8),
    to_signed(23, 8),
    to_signed(13, 8),
    to_signed(2, 8),
    to_signed(-8, 8),
    to_signed(-16, 8),
    to_signed(-16, 8),
    to_signed(-6, 8),
    to_signed(12, 8),
    to_signed(31, 8),
    to_signed(47, 8),
    to_signed(57, 8),
    to_signed(59, 8),
    to_signed(53, 8),
    to_signed(42, 8),
    to_signed(32, 8),
    to_signed(27, 8),
    to_signed(26, 8),
    to_signed(21, 8),
    to_signed(8, 8),
    to_signed(-15, 8),
    to_signed(-40, 8),
    to_signed(-60, 8),
    to_signed(-67, 8),
    to_signed(-58, 8),
    to_signed(-34, 8),
    to_signed(-7, 8),
    to_signed(13, 8),
    to_signed(17, 8),
    to_signed(8, 8),
    to_signed(-12, 8),
    to_signed(-35, 8),
    to_signed(-55, 8),
    to_signed(-68, 8),
    to_signed(-69, 8),
    to_signed(-56, 8),
    to_signed(-29, 8),
    to_signed(4, 8),
    to_signed(36, 8),
    to_signed(60, 8),
    to_signed(74, 8),
    to_signed(77, 8),
    to_signed(73, 8),
    to_signed(63, 8),
    to_signed(48, 8),
    to_signed(30, 8),
    to_signed(14, 8),
    to_signed(5, 8),
    to_signed(1, 8),
    to_signed(-2, 8),
    to_signed(-8, 8),
    to_signed(-19, 8),
    to_signed(-30, 8),
    to_signed(-37, 8),
    to_signed(-35, 8),
    to_signed(-28, 8),
    to_signed(-24, 8),
    to_signed(-26, 8),
    to_signed(-35, 8),
    to_signed(-46, 8),
    to_signed(-59, 8),
    to_signed(-67, 8),
    to_signed(-65, 8),
    to_signed(-51, 8),
    to_signed(-30, 8),
    to_signed(-10, 8),
    to_signed(6, 8),
    to_signed(17, 8),
    to_signed(23, 8),
    to_signed(23, 8),
    to_signed(18, 8),
    to_signed(13, 8),
    to_signed(13, 8),
    to_signed(20, 8),
    to_signed(29, 8),
    to_signed(35, 8),
    to_signed(34, 8),
    to_signed(28, 8),
    to_signed(18, 8),
    to_signed(6, 8),
    to_signed(-4, 8),
    to_signed(-12, 8),
    to_signed(-11, 8),
    to_signed(0, 8),
    to_signed(19, 8),
    to_signed(39, 8),
    to_signed(55, 8),
    to_signed(64, 8),
    to_signed(64, 8),
    to_signed(58, 8),
    to_signed(47, 8),
    to_signed(37, 8),
    to_signed(30, 8),
    to_signed(26, 8),
    to_signed(24, 8),
    to_signed(16, 8),
    to_signed(0, 8),
    to_signed(-24, 8),
    to_signed(-48, 8),
    to_signed(-62, 8),
    to_signed(-61, 8),
    to_signed(-43, 8),
    to_signed(-20, 8),
    to_signed(-2, 8),
    to_signed(3, 8),
    to_signed(-4, 8),
    to_signed(-22, 8),
    to_signed(-48, 8),
    to_signed(-75, 8),
    to_signed(-94, 8),
    to_signed(-97, 8),
    to_signed(-82, 8),
    to_signed(-53, 8),
    to_signed(-19, 8),
    to_signed(16, 8),
    to_signed(44, 8),
    to_signed(63, 8),
    to_signed(69, 8),
    to_signed(63, 8),
    to_signed(52, 8),
    to_signed(39, 8),
    to_signed(25, 8),
    to_signed(11, 8),
    to_signed(1, 8),
    to_signed(-4, 8),
    to_signed(-6, 8),
    to_signed(-10, 8),
    to_signed(-19, 8),
    to_signed(-32, 8),
    to_signed(-43, 8),
    to_signed(-44, 8),
    to_signed(-36, 8),
    to_signed(-28, 8),
    to_signed(-25, 8),
    to_signed(-29, 8),
    to_signed(-37, 8),
    to_signed(-48, 8),
    to_signed(-57, 8),
    to_signed(-58, 8),
    to_signed(-46, 8),
    to_signed(-25, 8),
    to_signed(0, 8),
    to_signed(22, 8),
    to_signed(37, 8),
    to_signed(44, 8),
    to_signed(44, 8),
    to_signed(38, 8),
    to_signed(30, 8),
    to_signed(26, 8),
    to_signed(27, 8),
    to_signed(31, 8),
    to_signed(33, 8),
    to_signed(31, 8),
    to_signed(24, 8),
    to_signed(13, 8),
    to_signed(2, 8),
    to_signed(-8, 8),
    to_signed(-16, 8),
    to_signed(-17, 8),
    to_signed(-9, 8),
    to_signed(9, 8),
    to_signed(29, 8),
    to_signed(46, 8),
    to_signed(57, 8),
    to_signed(61, 8),
    to_signed(59, 8),
    to_signed(50, 8),
    to_signed(38, 8),
    to_signed(28, 8),
    to_signed(22, 8),
    to_signed(19, 8),
    to_signed(12, 8),
    to_signed(-5, 8),
    to_signed(-31, 8),
    to_signed(-58, 8),
    to_signed(-73, 8),
    to_signed(-72, 8),
    to_signed(-53, 8),
    to_signed(-27, 8),
    to_signed(-3, 8),
    to_signed(8, 8),
    to_signed(4, 8),
    to_signed(-15, 8),
    to_signed(-41, 8),
    to_signed(-66, 8),
    to_signed(-80, 8),
    to_signed(-78, 8),
    to_signed(-61, 8),
    to_signed(-35, 8),
    to_signed(-4, 8),
    to_signed(27, 8),
    to_signed(53, 8),
    to_signed(71, 8),
    to_signed(77, 8),
    to_signed(74, 8),
    to_signed(66, 8),
    to_signed(55, 8),
    to_signed(41, 8),
    to_signed(23, 8),
    to_signed(8, 8),
    to_signed(0, 8),
    to_signed(-3, 8),
    to_signed(-6, 8),
    to_signed(-13, 8),
    to_signed(-23, 8),
    to_signed(-31, 8),
    to_signed(-32, 8),
    to_signed(-26, 8),
    to_signed(-18, 8),
    to_signed(-16, 8),
    to_signed(-22, 8),
    to_signed(-33, 8),
    to_signed(-47, 8),
    to_signed(-62, 8),
    to_signed(-69, 8),
    to_signed(-63, 8),
    to_signed(-45, 8),
    to_signed(-19, 8),
    to_signed(7, 8),
    to_signed(26, 8),
    to_signed(38, 8),
    to_signed(41, 8),
    to_signed(36, 8),
    to_signed(28, 8),
    to_signed(22, 8),
    to_signed(21, 8),
    to_signed(25, 8),
    to_signed(29, 8),
    to_signed(31, 8),
    to_signed(28, 8),
    to_signed(18, 8),
    to_signed(5, 8),
    to_signed(-7, 8),
    to_signed(-14, 8),
    to_signed(-12, 8),
    to_signed(-1, 8),
    to_signed(18, 8),
    to_signed(38, 8),
    to_signed(52, 8),
    to_signed(59, 8),
    to_signed(58, 8),
    to_signed(49, 8),
    to_signed(35, 8),
    to_signed(23, 8),
    to_signed(19, 8),
    to_signed(22, 8),
    to_signed(27, 8),
    to_signed(29, 8),
    to_signed(21, 8),
    to_signed(2, 8),
    to_signed(-26, 8),
    to_signed(-51, 8),
    to_signed(-64, 8),
    to_signed(-59, 8),
    to_signed(-40, 8),
    to_signed(-17, 8),
    to_signed(-3, 8),
    to_signed(-2, 8),
    to_signed(-14, 8),
    to_signed(-35, 8),
    to_signed(-59, 8),
    to_signed(-79, 8),
    to_signed(-88, 8),
    to_signed(-84, 8),
    to_signed(-66, 8),
    to_signed(-41, 8),
    to_signed(-14, 8),
    to_signed(11, 8),
    to_signed(34, 8),
    to_signed(49, 8),
    to_signed(56, 8),
    to_signed(55, 8),
    to_signed(50, 8),
    to_signed(40, 8),
    to_signed(25, 8),
    to_signed(7, 8),
    to_signed(-6, 8),
    to_signed(-13, 8),
    to_signed(-16, 8),
    to_signed(-17, 8),
    to_signed(-21, 8),
    to_signed(-26, 8),
    to_signed(-28, 8),
    to_signed(-23, 8),
    to_signed(-15, 8),
    to_signed(-13, 8),
    to_signed(-18, 8),
    to_signed(-28, 8),
    to_signed(-40, 8),
    to_signed(-51, 8),
    to_signed(-59, 8),
    to_signed(-56, 8),
    to_signed(-41, 8),
    to_signed(-16, 8),
    to_signed(10, 8),
    to_signed(32, 8),
    to_signed(46, 8),
    to_signed(51, 8),
    to_signed(48, 8),
    to_signed(38, 8),
    to_signed(28, 8),
    to_signed(22, 8),
    to_signed(23, 8),
    to_signed(27, 8),
    to_signed(31, 8),
    to_signed(30, 8),
    to_signed(22, 8),
    to_signed(9, 8),
    to_signed(-4, 8),
    to_signed(-13, 8),
    to_signed(-15, 8),
    to_signed(-10, 8),
    to_signed(4, 8),
    to_signed(23, 8),
    to_signed(40, 8),
    to_signed(52, 8),
    to_signed(57, 8),
    to_signed(54, 8),
    to_signed(44, 8),
    to_signed(32, 8),
    to_signed(23, 8),
    to_signed(19, 8),
    to_signed(18, 8),
    to_signed(18, 8),
    to_signed(12, 8),
    to_signed(-2, 8),
    to_signed(-27, 8),
    to_signed(-54, 8),
    to_signed(-72, 8),
    to_signed(-72, 8),
    to_signed(-56, 8),
    to_signed(-33, 8),
    to_signed(-14, 8),
    to_signed(-5, 8),
    to_signed(-9, 8),
    to_signed(-24, 8),
    to_signed(-44, 8),
    to_signed(-63, 8),
    to_signed(-74, 8),
    to_signed(-73, 8),
    to_signed(-57, 8),
    to_signed(-31, 8),
    to_signed(-1, 8),
    to_signed(29, 8),
    to_signed(55, 8),
    to_signed(73, 8),
    to_signed(79, 8),
    to_signed(77, 8),
    to_signed(68, 8),
    to_signed(56, 8),
    to_signed(41, 8),
    to_signed(24, 8),
    to_signed(11, 8),
    to_signed(4, 8),
    to_signed(1, 8),
    to_signed(-2, 8),
    to_signed(-9, 8),
    to_signed(-18, 8),
    to_signed(-24, 8),
    to_signed(-24, 8),
    to_signed(-18, 8),
    to_signed(-13, 8),
    to_signed(-14, 8),
    to_signed(-21, 8),
    to_signed(-33, 8),
    to_signed(-47, 8),
    to_signed(-58, 8),
    to_signed(-61, 8),
    to_signed(-53, 8),
    to_signed(-36, 8),
    to_signed(-15, 8),
    to_signed(6, 8),
    to_signed(25, 8),
    to_signed(38, 8),
    to_signed(43, 8),
    to_signed(40, 8),
    to_signed(32, 8),
    to_signed(26, 8),
    to_signed(23, 8),
    to_signed(24, 8),
    to_signed(27, 8),
    to_signed(30, 8),
    to_signed(29, 8),
    to_signed(21, 8),
    to_signed(9, 8),
    to_signed(-4, 8),
    to_signed(-13, 8),
    to_signed(-13, 8),
    to_signed(-4, 8),
    to_signed(11, 8),
    to_signed(27, 8),
    to_signed(41, 8),
    to_signed(50, 8),
    to_signed(52, 8),
    to_signed(44, 8),
    to_signed(30, 8),
    to_signed(19, 8),
    to_signed(14, 8),
    to_signed(15, 8),
    to_signed(16, 8),
    to_signed(16, 8),
    to_signed(11, 8),
    to_signed(-4, 8),
    to_signed(-26, 8),
    to_signed(-47, 8),
    to_signed(-57, 8),
    to_signed(-51, 8),
    to_signed(-35, 8),
    to_signed(-18, 8),
    to_signed(-9, 8),
    to_signed(-8, 8),
    to_signed(-15, 8),
    to_signed(-28, 8),
    to_signed(-44, 8),
    to_signed(-61, 8),
    to_signed(-71, 8),
    to_signed(-68, 8),
    to_signed(-51, 8),
    to_signed(-27, 8),
    to_signed(-1, 8),
    to_signed(25, 8),
    to_signed(48, 8),
    to_signed(63, 8),
    to_signed(66, 8),
    to_signed(61, 8),
    to_signed(51, 8),
    to_signed(38, 8),
    to_signed(23, 8),
    to_signed(8, 8),
    to_signed(-5, 8),
    to_signed(-13, 8),
    to_signed(-17, 8),
    to_signed(-20, 8),
    to_signed(-26, 8),
    to_signed(-32, 8),
    to_signed(-33, 8),
    to_signed(-26, 8),
    to_signed(-18, 8),
    to_signed(-15, 8),
    to_signed(-22, 8),
    to_signed(-34, 8),
    to_signed(-47, 8),
    to_signed(-59, 8),
    to_signed(-63, 8),
    to_signed(-57, 8),
    to_signed(-42, 8),
    to_signed(-20, 8),
    to_signed(5, 8),
    to_signed(27, 8),
    to_signed(43, 8),
    to_signed(50, 8),
    to_signed(48, 8),
    to_signed(40, 8),
    to_signed(31, 8),
    to_signed(24, 8),
    to_signed(22, 8),
    to_signed(25, 8),
    to_signed(31, 8),
    to_signed(35, 8),
    to_signed(32, 8),
    to_signed(23, 8),
    to_signed(9, 8),
    to_signed(-3, 8),
    to_signed(-9, 8),
    to_signed(-7, 8),
    to_signed(4, 8),
    to_signed(19, 8),
    to_signed(35, 8),
    to_signed(48, 8),
    to_signed(56, 8),
    to_signed(54, 8),
    to_signed(45, 8),
    to_signed(32, 8),
    to_signed(23, 8),
    to_signed(19, 8),
    to_signed(17, 8),
    to_signed(17, 8),
    to_signed(14, 8),
    to_signed(3, 8),
    to_signed(-18, 8),
    to_signed(-41, 8),
    to_signed(-56, 8),
    to_signed(-56, 8),
    to_signed(-43, 8),
    to_signed(-25, 8),
    to_signed(-9, 8),
    to_signed(-1, 8),
    to_signed(-3, 8),
    to_signed(-13, 8),
    to_signed(-30, 8),
    to_signed(-49, 8),
    to_signed(-65, 8),
    to_signed(-69, 8),
    to_signed(-58, 8),
    to_signed(-38, 8),
    to_signed(-12, 8),
    to_signed(14, 8),
    to_signed(37, 8),
    to_signed(52, 8),
    to_signed(56, 8),
    to_signed(51, 8),
    to_signed(43, 8),
    to_signed(33, 8),
    to_signed(22, 8),
    to_signed(12, 8),
    to_signed(3, 8),
    to_signed(-2, 8),
    to_signed(-5, 8),
    to_signed(-8, 8),
    to_signed(-15, 8),
    to_signed(-23, 8),
    to_signed(-26, 8),
    to_signed(-19, 8),
    to_signed(-7, 8),
    to_signed(1, 8),
    to_signed(0, 8),
    to_signed(-9, 8),
    to_signed(-24, 8),
    to_signed(-42, 8),
    to_signed(-55, 8),
    to_signed(-59, 8),
    to_signed(-52, 8),
    to_signed(-39, 8),
    to_signed(-21, 8),
    to_signed(-2, 8),
    to_signed(14, 8),
    to_signed(25, 8),
    to_signed(29, 8),
    to_signed(26, 8),
    to_signed(18, 8),
    to_signed(10, 8),
    to_signed(6, 8),
    to_signed(9, 8),
    to_signed(15, 8),
    to_signed(23, 8),
    to_signed(27, 8),
    to_signed(24, 8),
    to_signed(14, 8),
    to_signed(1, 8),
    to_signed(-8, 8),
    to_signed(-9, 8),
    to_signed(0, 8),
    to_signed(15, 8),
    to_signed(32, 8),
    to_signed(46, 8),
    to_signed(54, 8),
    to_signed(54, 8),
    to_signed(45, 8),
    to_signed(31, 8),
    to_signed(19, 8),
    to_signed(14, 8),
    to_signed(15, 8),
    to_signed(17, 8),
    to_signed(15, 8),
    to_signed(7, 8),
    to_signed(-11, 8),
    to_signed(-37, 8),
    to_signed(-60, 8),
    to_signed(-69, 8),
    to_signed(-63, 8),
    to_signed(-45, 8),
    to_signed(-25, 8),
    to_signed(-9, 8),
    to_signed(-2, 8),
    to_signed(-7, 8),
    to_signed(-20, 8),
    to_signed(-39, 8),
    to_signed(-59, 8),
    to_signed(-73, 8),
    to_signed(-72, 8),
    to_signed(-55, 8),
    to_signed(-28, 8),
    to_signed(3, 8),
    to_signed(33, 8),
    to_signed(56, 8),
    to_signed(68, 8),
    to_signed(67, 8),
    to_signed(59, 8),
    to_signed(47, 8),
    to_signed(35, 8),
    to_signed(24, 8),
    to_signed(14, 8),
    to_signed(5, 8),
    to_signed(-2, 8),
    to_signed(-6, 8),
    to_signed(-11, 8),
    to_signed(-17, 8),
    to_signed(-23, 8),
    to_signed(-23, 8),
    to_signed(-18, 8),
    to_signed(-11, 8),
    to_signed(-10, 8),
    to_signed(-14, 8),
    to_signed(-24, 8),
    to_signed(-36, 8),
    to_signed(-46, 8),
    to_signed(-50, 8),
    to_signed(-46, 8),
    to_signed(-36, 8),
    to_signed(-20, 8),
    to_signed(-2, 8),
    to_signed(17, 8),
    to_signed(30, 8),
    to_signed(35, 8),
    to_signed(34, 8),
    to_signed(26, 8),
    to_signed(16, 8),
    to_signed(9, 8),
    to_signed(10, 8),
    to_signed(17, 8),
    to_signed(26, 8),
    to_signed(31, 8),
    to_signed(29, 8),
    to_signed(17, 8),
    to_signed(0, 8),
    to_signed(-17, 8),
    to_signed(-27, 8),
    to_signed(-24, 8),
    to_signed(-10, 8),
    to_signed(13, 8),
    to_signed(36, 8),
    to_signed(53, 8),
    to_signed(59, 8),
    to_signed(56, 8),
    to_signed(45, 8),
    to_signed(33, 8),
    to_signed(25, 8),
    to_signed(24, 8),
    to_signed(27, 8),
    to_signed(29, 8),
    to_signed(27, 8),
    to_signed(17, 8),
    to_signed(-2, 8),
    to_signed(-27, 8),
    to_signed(-45, 8),
    to_signed(-50, 8),
    to_signed(-39, 8),
    to_signed(-20, 8),
    to_signed(1, 8),
    to_signed(14, 8),
    to_signed(14, 8),
    to_signed(2, 8),
    to_signed(-17, 8),
    to_signed(-38, 8),
    to_signed(-57, 8),
    to_signed(-65, 8),
    to_signed(-59, 8),
    to_signed(-39, 8),
    to_signed(-12, 8),
    to_signed(15, 8),
    to_signed(38, 8),
    to_signed(53, 8),
    to_signed(57, 8),
    to_signed(51, 8),
    to_signed(40, 8),
    to_signed(29, 8),
    to_signed(19, 8),
    to_signed(10, 8),
    to_signed(3, 8),
    to_signed(-3, 8),
    to_signed(-9, 8),
    to_signed(-15, 8),
    to_signed(-22, 8),
    to_signed(-30, 8),
    to_signed(-36, 8),
    to_signed(-35, 8),
    to_signed(-29, 8),
    to_signed(-23, 8),
    to_signed(-23, 8),
    to_signed(-29, 8),
    to_signed(-41, 8),
    to_signed(-56, 8),
    to_signed(-70, 8),
    to_signed(-74, 8),
    to_signed(-69, 8),
    to_signed(-55, 8),
    to_signed(-36, 8),
    to_signed(-12, 8),
    to_signed(8, 8),
    to_signed(22, 8),
    to_signed(27, 8),
    to_signed(25, 8),
    to_signed(19, 8),
    to_signed(13, 8),
    to_signed(11, 8),
    to_signed(16, 8),
    to_signed(24, 8),
    to_signed(31, 8),
    to_signed(35, 8),
    to_signed(36, 8),
    to_signed(28, 8),
    to_signed(13, 8),
    to_signed(-1, 8),
    to_signed(-9, 8),
    to_signed(-4, 8),
    to_signed(10, 8),
    to_signed(31, 8),
    to_signed(50, 8),
    to_signed(61, 8),
    to_signed(63, 8),
    to_signed(56, 8),
    to_signed(44, 8),
    to_signed(34, 8),
    to_signed(30, 8),
    to_signed(34, 8),
    to_signed(40, 8),
    to_signed(46, 8),
    to_signed(46, 8),
    to_signed(35, 8),
    to_signed(10, 8),
    to_signed(-20, 8),
    to_signed(-45, 8),
    to_signed(-54, 8),
    to_signed(-47, 8),
    to_signed(-28, 8),
    to_signed(-8, 8),
    to_signed(6, 8),
    to_signed(8, 8),
    to_signed(-2, 8),
    to_signed(-23, 8),
    to_signed(-49, 8),
    to_signed(-74, 8),
    to_signed(-86, 8),
    to_signed(-83, 8),
    to_signed(-66, 8),
    to_signed(-43, 8),
    to_signed(-17, 8),
    to_signed(8, 8),
    to_signed(25, 8),
    to_signed(33, 8),
    to_signed(30, 8),
    to_signed(24, 8),
    to_signed(18, 8),
    to_signed(12, 8),
    to_signed(6, 8),
    to_signed(0, 8),
    to_signed(-8, 8),
    to_signed(-15, 8),
    to_signed(-21, 8),
    to_signed(-26, 8),
    to_signed(-30, 8),
    to_signed(-32, 8),
    to_signed(-28, 8),
    to_signed(-21, 8),
    to_signed(-14, 8),
    to_signed(-12, 8),
    to_signed(-15, 8),
    to_signed(-23, 8),
    to_signed(-34, 8),
    to_signed(-42, 8),
    to_signed(-44, 8),
    to_signed(-40, 8),
    to_signed(-29, 8),
    to_signed(-11, 8),
    to_signed(9, 8),
    to_signed(25, 8),
    to_signed(35, 8),
    to_signed(40, 8),
    to_signed(40, 8),
    to_signed(37, 8),
    to_signed(33, 8),
    to_signed(32, 8),
    to_signed(35, 8),
    to_signed(39, 8),
    to_signed(42, 8),
    to_signed(42, 8),
    to_signed(37, 8),
    to_signed(26, 8),
    to_signed(12, 8),
    to_signed(0, 8),
    to_signed(-6, 8),
    to_signed(-3, 8),
    to_signed(11, 8),
    to_signed(30, 8),
    to_signed(49, 8),
    to_signed(59, 8),
    to_signed(60, 8),
    to_signed(51, 8),
    to_signed(38, 8),
    to_signed(25, 8),
    to_signed(17, 8),
    to_signed(13, 8),
    to_signed(12, 8),
    to_signed(12, 8),
    to_signed(6, 8),
    to_signed(-10, 8),
    to_signed(-36, 8),
    to_signed(-63, 8),
    to_signed(-79, 8),
    to_signed(-79, 8),
    to_signed(-62, 8),
    to_signed(-35, 8),
    to_signed(-10, 8),
    to_signed(3, 8),
    to_signed(0, 8),
    to_signed(-17, 8),
    to_signed(-40, 8),
    to_signed(-63, 8),
    to_signed(-78, 8),
    to_signed(-79, 8),
    to_signed(-65, 8),
    to_signed(-40, 8),
    to_signed(-10, 8),
    to_signed(18, 8),
    to_signed(40, 8),
    to_signed(54, 8),
    to_signed(57, 8),
    to_signed(52, 8),
    to_signed(45, 8),
    to_signed(36, 8),
    to_signed(26, 8),
    to_signed(17, 8),
    to_signed(8, 8),
    to_signed(1, 8),
    to_signed(-4, 8),
    to_signed(-8, 8),
    to_signed(-13, 8),
    to_signed(-19, 8),
    to_signed(-21, 8),
    to_signed(-17, 8),
    to_signed(-8, 8),
    to_signed(-1, 8),
    to_signed(0, 8),
    to_signed(-7, 8),
    to_signed(-20, 8),
    to_signed(-35, 8),
    to_signed(-48, 8),
    to_signed(-54, 8),
    to_signed(-51, 8),
    to_signed(-39, 8),
    to_signed(-19, 8),
    to_signed(1, 8),
    to_signed(16, 8),
    to_signed(24, 8),
    to_signed(26, 8),
    to_signed(23, 8),
    to_signed(19, 8),
    to_signed(16, 8),
    to_signed(17, 8),
    to_signed(20, 8),
    to_signed(22, 8),
    to_signed(21, 8),
    to_signed(17, 8),
    to_signed(11, 8),
    to_signed(1, 8),
    to_signed(-10, 8),
    to_signed(-19, 8),
    to_signed(-20, 8),
    to_signed(-11, 8),
    to_signed(8, 8),
    to_signed(29, 8),
    to_signed(45, 8),
    to_signed(54, 8),
    to_signed(53, 8),
    to_signed(44, 8),
    to_signed(31, 8),
    to_signed(19, 8),
    to_signed(11, 8),
    to_signed(9, 8),
    to_signed(11, 8),
    to_signed(12, 8),
    to_signed(6, 8),
    to_signed(-11, 8),
    to_signed(-35, 8),
    to_signed(-58, 8),
    to_signed(-69, 8),
    to_signed(-61, 8),
    to_signed(-40, 8),
    to_signed(-16, 8),
    to_signed(0, 8),
    to_signed(2, 8),
    to_signed(-7, 8),
    to_signed(-27, 8),
    to_signed(-52, 8),
    to_signed(-72, 8),
    to_signed(-81, 8),
    to_signed(-74, 8),
    to_signed(-52, 8),
    to_signed(-23, 8),
    to_signed(7, 8),
    to_signed(33, 8),
    to_signed(51, 8),
    to_signed(59, 8),
    to_signed(55, 8),
    to_signed(45, 8),
    to_signed(33, 8),
    to_signed(21, 8),
    to_signed(9, 8),
    to_signed(-2, 8),
    to_signed(-11, 8),
    to_signed(-17, 8),
    to_signed(-21, 8),
    to_signed(-26, 8),
    to_signed(-34, 8),
    to_signed(-42, 8),
    to_signed(-43, 8),
    to_signed(-37, 8),
    to_signed(-29, 8),
    to_signed(-24, 8),
    to_signed(-26, 8),
    to_signed(-34, 8),
    to_signed(-46, 8),
    to_signed(-59, 8),
    to_signed(-67, 8),
    to_signed(-64, 8),
    to_signed(-49, 8),
    to_signed(-26, 8),
    to_signed(-1, 8),
    to_signed(19, 8),
    to_signed(32, 8),
    to_signed(37, 8),
    to_signed(34, 8),
    to_signed(26, 8),
    to_signed(19, 8),
    to_signed(18, 8),
    to_signed(23, 8),
    to_signed(30, 8),
    to_signed(34, 8),
    to_signed(32, 8),
    to_signed(25, 8),
    to_signed(15, 8),
    to_signed(4, 8),
    to_signed(-7, 8),
    to_signed(-12, 8),
    to_signed(-9, 8),
    to_signed(4, 8),
    to_signed(24, 8),
    to_signed(45, 8),
    to_signed(62, 8),
    to_signed(69, 8),
    to_signed(67, 8),
    to_signed(57, 8),
    to_signed(44, 8),
    to_signed(32, 8),
    to_signed(26, 8),
    to_signed(25, 8),
    to_signed(29, 8),
    to_signed(29, 8),
    to_signed(19, 8),
    to_signed(-4, 8),
    to_signed(-34, 8),
    to_signed(-59, 8),
    to_signed(-67, 8),
    to_signed(-56, 8),
    to_signed(-34, 8),
    to_signed(-13, 8),
    to_signed(0, 8),
    to_signed(0, 8),
    to_signed(-12, 8),
    to_signed(-33, 8),
    to_signed(-56, 8),
    to_signed(-73, 8),
    to_signed(-79, 8),
    to_signed(-70, 8),
    to_signed(-48, 8),
    to_signed(-20, 8),
    to_signed(8, 8),
    to_signed(30, 8),
    to_signed(44, 8),
    to_signed(47, 8),
    to_signed(44, 8),
    to_signed(37, 8),
    to_signed(27, 8),
    to_signed(15, 8),
    to_signed(2, 8),
    to_signed(-9, 8),
    to_signed(-15, 8),
    to_signed(-18, 8),
    to_signed(-19, 8),
    to_signed(-23, 8),
    to_signed(-29, 8),
    to_signed(-34, 8),
    to_signed(-32, 8),
    to_signed(-23, 8),
    to_signed(-14, 8),
    to_signed(-9, 8),
    to_signed(-13, 8),
    to_signed(-24, 8),
    to_signed(-39, 8),
    to_signed(-51, 8),
    to_signed(-55, 8),
    to_signed(-50, 8),
    to_signed(-36, 8),
    to_signed(-16, 8),
    to_signed(6, 8),
    to_signed(26, 8),
    to_signed(38, 8),
    to_signed(40, 8),
    to_signed(35, 8),
    to_signed(26, 8),
    to_signed(20, 8),
    to_signed(20, 8),
    to_signed(25, 8),
    to_signed(31, 8),
    to_signed(34, 8),
    to_signed(33, 8),
    to_signed(27, 8),
    to_signed(18, 8),
    to_signed(7, 8),
    to_signed(-1, 8),
    to_signed(-4, 8),
    to_signed(1, 8),
    to_signed(13, 8),
    to_signed(30, 8),
    to_signed(45, 8),
    to_signed(55, 8),
    to_signed(58, 8),
    to_signed(53, 8),
    to_signed(43, 8),
    to_signed(29, 8),
    to_signed(17, 8),
    to_signed(12, 8),
    to_signed(14, 8),
    to_signed(18, 8),
    to_signed(16, 8),
    to_signed(0, 8),
    to_signed(-28, 8),
    to_signed(-56, 8),
    to_signed(-74, 8),
    to_signed(-72, 8),
    to_signed(-56, 8),
    to_signed(-33, 8),
    to_signed(-14, 8),
    to_signed(-3, 8),
    to_signed(-3, 8),
    to_signed(-15, 8),
    to_signed(-34, 8),
    to_signed(-55, 8),
    to_signed(-70, 8),
    to_signed(-74, 8),
    to_signed(-62, 8),
    to_signed(-38, 8),
    to_signed(-7, 8),
    to_signed(22, 8),
    to_signed(46, 8),
    to_signed(59, 8),
    to_signed(63, 8),
    to_signed(60, 8),
    to_signed(51, 8),
    to_signed(38, 8),
    to_signed(21, 8),
    to_signed(5, 8),
    to_signed(-6, 8),
    to_signed(-11, 8),
    to_signed(-12, 8),
    to_signed(-12, 8),
    to_signed(-17, 8),
    to_signed(-23, 8),
    to_signed(-25, 8),
    to_signed(-20, 8),
    to_signed(-14, 8),
    to_signed(-13, 8),
    to_signed(-16, 8),
    to_signed(-24, 8),
    to_signed(-34, 8),
    to_signed(-44, 8),
    to_signed(-49, 8),
    to_signed(-46, 8),
    to_signed(-33, 8),
    to_signed(-14, 8),
    to_signed(7, 8),
    to_signed(24, 8),
    to_signed(36, 8),
    to_signed(41, 8),
    to_signed(40, 8),
    to_signed(35, 8),
    to_signed(28, 8),
    to_signed(25, 8),
    to_signed(31, 8),
    to_signed(40, 8),
    to_signed(46, 8),
    to_signed(44, 8),
    to_signed(35, 8),
    to_signed(20, 8),
    to_signed(5, 8),
    to_signed(-6, 8),
    to_signed(-10, 8),
    to_signed(-6, 8),
    to_signed(7, 8),
    to_signed(26, 8),
    to_signed(47, 8),
    to_signed(62, 8),
    to_signed(70, 8),
    to_signed(71, 8),
    to_signed(64, 8),
    to_signed(51, 8),
    to_signed(37, 8),
    to_signed(27, 8),
    to_signed(23, 8),
    to_signed(24, 8),
    to_signed(23, 8),
    to_signed(14, 8),
    to_signed(-6, 8),
    to_signed(-31, 8),
    to_signed(-49, 8),
    to_signed(-53, 8),
    to_signed(-42, 8),
    to_signed(-24, 8),
    to_signed(-7, 8),
    to_signed(3, 8),
    to_signed(2, 8),
    to_signed(-9, 8),
    to_signed(-28, 8),
    to_signed(-48, 8),
    to_signed(-64, 8),
    to_signed(-69, 8),
    to_signed(-58, 8),
    to_signed(-35, 8),
    to_signed(-6, 8),
    to_signed(23, 8),
    to_signed(48, 8),
    to_signed(64, 8),
    to_signed(67, 8),
    to_signed(62, 8),
    to_signed(53, 8),
    to_signed(39, 8),
    to_signed(22, 8),
    to_signed(6, 8),
    to_signed(-8, 8),
    to_signed(-16, 8),
    to_signed(-18, 8),
    to_signed(-16, 8),
    to_signed(-16, 8),
    to_signed(-21, 8),
    to_signed(-25, 8),
    to_signed(-22, 8),
    to_signed(-15, 8),
    to_signed(-11, 8),
    to_signed(-14, 8),
    to_signed(-22, 8),
    to_signed(-34, 8),
    to_signed(-46, 8),
    to_signed(-54, 8),
    to_signed(-53, 8),
    to_signed(-43, 8),
    to_signed(-25, 8),
    to_signed(-3, 8),
    to_signed(20, 8),
    to_signed(37, 8),
    to_signed(46, 8),
    to_signed(45, 8),
    to_signed(38, 8),
    to_signed(27, 8),
    to_signed(18, 8),
    to_signed(19, 8),
    to_signed(29, 8),
    to_signed(40, 8),
    to_signed(46, 8),
    to_signed(44, 8),
    to_signed(34, 8),
    to_signed(18, 8),
    to_signed(3, 8),
    to_signed(-8, 8),
    to_signed(-11, 8),
    to_signed(-6, 8),
    to_signed(9, 8),
    to_signed(29, 8),
    to_signed(47, 8),
    to_signed(57, 8),
    to_signed(59, 8),
    to_signed(53, 8),
    to_signed(40, 8),
    to_signed(23, 8),
    to_signed(9, 8),
    to_signed(4, 8),
    to_signed(5, 8),
    to_signed(9, 8),
    to_signed(7, 8),
    to_signed(-6, 8),
    to_signed(-30, 8),
    to_signed(-53, 8),
    to_signed(-64, 8),
    to_signed(-59, 8),
    to_signed(-45, 8),
    to_signed(-26, 8),
    to_signed(-10, 8),
    to_signed(-1, 8),
    to_signed(-5, 8),
    to_signed(-18, 8),
    to_signed(-38, 8),
    to_signed(-59, 8),
    to_signed(-73, 8),
    to_signed(-74, 8),
    to_signed(-61, 8),
    to_signed(-36, 8),
    to_signed(-5, 8),
    to_signed(25, 8),
    to_signed(49, 8),
    to_signed(60, 8),
    to_signed(61, 8),
    to_signed(56, 8),
    to_signed(45, 8),
    to_signed(29, 8),
    to_signed(9, 8),
    to_signed(-6, 8),
    to_signed(-14, 8),
    to_signed(-16, 8),
    to_signed(-16, 8),
    to_signed(-18, 8),
    to_signed(-24, 8),
    to_signed(-29, 8),
    to_signed(-28, 8),
    to_signed(-21, 8),
    to_signed(-15, 8),
    to_signed(-15, 8),
    to_signed(-21, 8),
    to_signed(-32, 8),
    to_signed(-45, 8),
    to_signed(-58, 8),
    to_signed(-64, 8),
    to_signed(-60, 8),
    to_signed(-45, 8),
    to_signed(-22, 8),
    to_signed(4, 8),
    to_signed(28, 8),
    to_signed(43, 8),
    to_signed(49, 8),
    to_signed(46, 8),
    to_signed(35, 8),
    to_signed(20, 8),
    to_signed(9, 8),
    to_signed(10, 8),
    to_signed(18, 8),
    to_signed(26, 8),
    to_signed(29, 8),
    to_signed(24, 8),
    to_signed(13, 8),
    to_signed(-2, 8),
    to_signed(-14, 8),
    to_signed(-19, 8),
    to_signed(-17, 8),
    to_signed(-6, 8),
    to_signed(15, 8),
    to_signed(39, 8),
    to_signed(58, 8),
    to_signed(68, 8),
    to_signed(68, 8),
    to_signed(59, 8),
    to_signed(44, 8),
    to_signed(30, 8),
    to_signed(24, 8),
    to_signed(27, 8),
    to_signed(34, 8),
    to_signed(37, 8),
    to_signed(29, 8),
    to_signed(8, 8),
    to_signed(-21, 8),
    to_signed(-43, 8),
    to_signed(-51, 8),
    to_signed(-46, 8),
    to_signed(-32, 8),
    to_signed(-17, 8),
    to_signed(-4, 8),
    to_signed(0, 8),
    to_signed(-7, 8),
    to_signed(-25, 8),
    to_signed(-46, 8),
    to_signed(-65, 8),
    to_signed(-75, 8),
    to_signed(-70, 8),
    to_signed(-52, 8),
    to_signed(-26, 8),
    to_signed(4, 8),
    to_signed(32, 8),
    to_signed(51, 8),
    to_signed(59, 8),
    to_signed(56, 8),
    to_signed(45, 8),
    to_signed(30, 8),
    to_signed(10, 8),
    to_signed(-8, 8),
    to_signed(-21, 8),
    to_signed(-27, 8),
    to_signed(-29, 8),
    to_signed(-31, 8),
    to_signed(-36, 8),
    to_signed(-43, 8),
    to_signed(-46, 8),
    to_signed(-41, 8),
    to_signed(-31, 8),
    to_signed(-23, 8),
    to_signed(-23, 8),
    to_signed(-29, 8),
    to_signed(-39, 8),
    to_signed(-50, 8),
    to_signed(-58, 8),
    to_signed(-57, 8),
    to_signed(-46, 8),
    to_signed(-28, 8),
    to_signed(-5, 8),
    to_signed(18, 8),
    to_signed(36, 8),
    to_signed(46, 8),
    to_signed(47, 8),
    to_signed(41, 8),
    to_signed(30, 8),
    to_signed(20, 8),
    to_signed(18, 8),
    to_signed(24, 8),
    to_signed(34, 8),
    to_signed(39, 8),
    to_signed(38, 8),
    to_signed(30, 8),
    to_signed(18, 8),
    to_signed(5, 8),
    to_signed(-4, 8),
    to_signed(-6, 8),
    to_signed(-1, 8),
    to_signed(13, 8),
    to_signed(34, 8),
    to_signed(55, 8),
    to_signed(68, 8),
    to_signed(70, 8),
    to_signed(62, 8),
    to_signed(46, 8),
    to_signed(28, 8),
    to_signed(16, 8),
    to_signed(11, 8),
    to_signed(12, 8),
    to_signed(13, 8),
    to_signed(6, 8),
    to_signed(-13, 8),
    to_signed(-41, 8),
    to_signed(-64, 8),
    to_signed(-75, 8),
    to_signed(-69, 8),
    to_signed(-52, 8),
    to_signed(-30, 8),
    to_signed(-13, 8),
    to_signed(-8, 8),
    to_signed(-16, 8),
    to_signed(-35, 8),
    to_signed(-59, 8),
    to_signed(-81, 8),
    to_signed(-95, 8),
    to_signed(-95, 8),
    to_signed(-80, 8),
    to_signed(-55, 8),
    to_signed(-24, 8),
    to_signed(5, 8),
    to_signed(27, 8),
    to_signed(40, 8),
    to_signed(43, 8),
    to_signed(39, 8),
    to_signed(30, 8),
    to_signed(15, 8),
    to_signed(0, 8),
    to_signed(-11, 8),
    to_signed(-15, 8),
    to_signed(-14, 8),
    to_signed(-12, 8),
    to_signed(-15, 8),
    to_signed(-19, 8),
    to_signed(-20, 8),
    to_signed(-14, 8),
    to_signed(-2, 8),
    to_signed(7, 8),
    to_signed(10, 8),
    to_signed(3, 8),
    to_signed(-11, 8),
    to_signed(-28, 8),
    to_signed(-43, 8),
    to_signed(-48, 8),
    to_signed(-43, 8),
    to_signed(-28, 8),
    to_signed(-6, 8),
    to_signed(16, 8),
    to_signed(33, 8),
    to_signed(42, 8),
    to_signed(42, 8),
    to_signed(34, 8),
    to_signed(21, 8),
    to_signed(7, 8),
    to_signed(-1, 8),
    to_signed(2, 8),
    to_signed(10, 8),
    to_signed(17, 8),
    to_signed(20, 8),
    to_signed(16, 8),
    to_signed(6, 8),
    to_signed(-6, 8),
    to_signed(-16, 8),
    to_signed(-20, 8),
    to_signed(-17, 8),
    to_signed(-7, 8),
    to_signed(12, 8),
    to_signed(35, 8),
    to_signed(54, 8),
    to_signed(64, 8),
    to_signed(61, 8),
    to_signed(48, 8),
    to_signed(32, 8),
    to_signed(18, 8),
    to_signed(12, 8),
    to_signed(12, 8),
    to_signed(15, 8),
    to_signed(14, 8),
    to_signed(2, 8),
    to_signed(-22, 8),
    to_signed(-49, 8),
    to_signed(-67, 8),
    to_signed(-69, 8),
    to_signed(-56, 8),
    to_signed(-36, 8),
    to_signed(-16, 8),
    to_signed(-4, 8),
    to_signed(-4, 8),
    to_signed(-15, 8),
    to_signed(-33, 8),
    to_signed(-54, 8),
    to_signed(-68, 8),
    to_signed(-70, 8),
    to_signed(-57, 8),
    to_signed(-35, 8),
    to_signed(-10, 8),
    to_signed(15, 8),
    to_signed(38, 8),
    to_signed(54, 8),
    to_signed(61, 8),
    to_signed(60, 8),
    to_signed(54, 8),
    to_signed(43, 8),
    to_signed(29, 8),
    to_signed(14, 8),
    to_signed(2, 8),
    to_signed(-5, 8),
    to_signed(-9, 8),
    to_signed(-15, 8),
    to_signed(-25, 8),
    to_signed(-32, 8),
    to_signed(-32, 8),
    to_signed(-22, 8),
    to_signed(-8, 8),
    to_signed(3, 8),
    to_signed(5, 8),
    to_signed(-4, 8),
    to_signed(-21, 8),
    to_signed(-39, 8),
    to_signed(-51, 8),
    to_signed(-52, 8),
    to_signed(-41, 8),
    to_signed(-23, 8),
    to_signed(-1, 8),
    to_signed(18, 8),
    to_signed(30, 8),
    to_signed(34, 8),
    to_signed(31, 8),
    to_signed(20, 8),
    to_signed(8, 8),
    to_signed(0, 8),
    to_signed(2, 8),
    to_signed(12, 8),
    to_signed(24, 8),
    to_signed(31, 8),
    to_signed(32, 8),
    to_signed(26, 8),
    to_signed(16, 8),
    to_signed(5, 8),
    to_signed(-2, 8),
    to_signed(-4, 8),
    to_signed(2, 8),
    to_signed(15, 8),
    to_signed(35, 8),
    to_signed(57, 8),
    to_signed(73, 8),
    to_signed(78, 8),
    to_signed(71, 8),
    to_signed(56, 8),
    to_signed(41, 8),
    to_signed(31, 8),
    to_signed(27, 8),
    to_signed(27, 8),
    to_signed(24, 8),
    to_signed(14, 8),
    to_signed(-7, 8),
    to_signed(-34, 8),
    to_signed(-59, 8),
    to_signed(-70, 8),
    to_signed(-63, 8),
    to_signed(-43, 8),
    to_signed(-19, 8),
    to_signed(0, 8),
    to_signed(7, 8),
    to_signed(0, 8),
    to_signed(-18, 8),
    to_signed(-41, 8),
    to_signed(-62, 8),
    to_signed(-74, 8),
    to_signed(-71, 8),
    to_signed(-54, 8),
    to_signed(-30, 8),
    to_signed(-2, 8),
    to_signed(24, 8),
    to_signed(45, 8),
    to_signed(56, 8),
    to_signed(58, 8),
    to_signed(52, 8),
    to_signed(39, 8),
    to_signed(21, 8),
    to_signed(2, 8),
    to_signed(-12, 8),
    to_signed(-17, 8),
    to_signed(-16, 8),
    to_signed(-14, 8),
    to_signed(-17, 8),
    to_signed(-23, 8),
    to_signed(-27, 8),
    to_signed(-24, 8),
    to_signed(-15, 8),
    to_signed(-6, 8),
    to_signed(-2, 8),
    to_signed(-6, 8),
    to_signed(-19, 8),
    to_signed(-35, 8),
    to_signed(-49, 8),
    to_signed(-53, 8),
    to_signed(-44, 8),
    to_signed(-25, 8),
    to_signed(-2, 8),
    to_signed(19, 8),
    to_signed(34, 8),
    to_signed(41, 8),
    to_signed(40, 8),
    to_signed(30, 8),
    to_signed(17, 8),
    to_signed(6, 8),
    to_signed(4, 8),
    to_signed(11, 8),
    to_signed(23, 8),
    to_signed(33, 8),
    to_signed(38, 8),
    to_signed(36, 8),
    to_signed(27, 8),
    to_signed(14, 8),
    to_signed(1, 8),
    to_signed(-8, 8),
    to_signed(-9, 8),
    to_signed(-3, 8),
    to_signed(11, 8),
    to_signed(29, 8),
    to_signed(46, 8),
    to_signed(56, 8),
    to_signed(55, 8),
    to_signed(45, 8),
    to_signed(31, 8),
    to_signed(20, 8),
    to_signed(16, 8),
    to_signed(17, 8),
    to_signed(19, 8),
    to_signed(15, 8),
    to_signed(1, 8),
    to_signed(-24, 8),
    to_signed(-52, 8),
    to_signed(-74, 8),
    to_signed(-80, 8),
    to_signed(-68, 8),
    to_signed(-45, 8),
    to_signed(-20, 8),
    to_signed(-3, 8),
    to_signed(4, 8),
    to_signed(-3, 8),
    to_signed(-20, 8),
    to_signed(-43, 8),
    to_signed(-62, 8),
    to_signed(-70, 8),
    to_signed(-64, 8),
    to_signed(-49, 8),
    to_signed(-30, 8),
    to_signed(-8, 8),
    to_signed(15, 8),
    to_signed(36, 8),
    to_signed(48, 8),
    to_signed(51, 8),
    to_signed(46, 8),
    to_signed(33, 8),
    to_signed(17, 8),
    to_signed(2, 8),
    to_signed(-8, 8),
    to_signed(-12, 8),
    to_signed(-13, 8),
    to_signed(-14, 8),
    to_signed(-19, 8),
    to_signed(-25, 8),
    to_signed(-28, 8),
    to_signed(-20, 8),
    to_signed(-6, 8),
    to_signed(7, 8),
    to_signed(12, 8),
    to_signed(6, 8),
    to_signed(-9, 8),
    to_signed(-28, 8),
    to_signed(-44, 8),
    to_signed(-49, 8),
    to_signed(-40, 8),
    to_signed(-23, 8),
    to_signed(-2, 8),
    to_signed(16, 8),
    to_signed(27, 8),
    to_signed(30, 8),
    to_signed(25, 8),
    to_signed(15, 8),
    to_signed(2, 8),
    to_signed(-6, 8),
    to_signed(-6, 8),
    to_signed(2, 8),
    to_signed(14, 8),
    to_signed(25, 8),
    to_signed(31, 8),
    to_signed(31, 8),
    to_signed(24, 8),
    to_signed(15, 8),
    to_signed(8, 8),
    to_signed(4, 8),
    to_signed(7, 8),
    to_signed(16, 8),
    to_signed(32, 8),
    to_signed(50, 8),
    to_signed(62, 8),
    to_signed(66, 8),
    to_signed(60, 8),
    to_signed(46, 8),
    to_signed(32, 8),
    to_signed(26, 8),
    to_signed(28, 8),
    to_signed(35, 8),
    to_signed(39, 8),
    to_signed(35, 8),
    to_signed(18, 8),
    to_signed(-10, 8),
    to_signed(-42, 8),
    to_signed(-66, 8),
    to_signed(-73, 8),
    to_signed(-61, 8),
    to_signed(-38, 8),
    to_signed(-12, 8),
    to_signed(9, 8),
    to_signed(18, 8),
    to_signed(12, 8),
    to_signed(-6, 8),
    to_signed(-30, 8),
    to_signed(-50, 8),
    to_signed(-59, 8),
    to_signed(-57, 8),
    to_signed(-46, 8),
    to_signed(-27, 8),
    to_signed(-5, 8),
    to_signed(18, 8),
    to_signed(35, 8),
    to_signed(44, 8),
    to_signed(44, 8),
    to_signed(36, 8),
    to_signed(23, 8),
    to_signed(9, 8),
    to_signed(-3, 8),
    to_signed(-10, 8),
    to_signed(-13, 8),
    to_signed(-14, 8),
    to_signed(-18, 8),
    to_signed(-26, 8),
    to_signed(-33, 8),
    to_signed(-34, 8),
    to_signed(-23, 8),
    to_signed(-7, 8),
    to_signed(7, 8),
    to_signed(11, 8),
    to_signed(3, 8),
    to_signed(-15, 8),
    to_signed(-37, 8),
    to_signed(-55, 8),
    to_signed(-59, 8),
    to_signed(-51, 8),
    to_signed(-33, 8),
    to_signed(-12, 8),
    to_signed(5, 8),
    to_signed(16, 8),
    to_signed(18, 8),
    to_signed(12, 8),
    to_signed(2, 8),
    to_signed(-8, 8),
    to_signed(-13, 8),
    to_signed(-9, 8),
    to_signed(2, 8),
    to_signed(16, 8),
    to_signed(26, 8),
    to_signed(28, 8),
    to_signed(24, 8),
    to_signed(15, 8),
    to_signed(6, 8),
    to_signed(0, 8),
    to_signed(1, 8),
    to_signed(11, 8),
    to_signed(28, 8),
    to_signed(47, 8),
    to_signed(63, 8),
    to_signed(70, 8),
    to_signed(66, 8),
    to_signed(53, 8),
    to_signed(36, 8),
    to_signed(23, 8),
    to_signed(19, 8),
    to_signed(26, 8),
    to_signed(38, 8),
    to_signed(46, 8),
    to_signed(45, 8),
    to_signed(28, 8),
    to_signed(-4, 8),
    to_signed(-43, 8),
    to_signed(-74, 8),
    to_signed(-87, 8),
    to_signed(-81, 8),
    to_signed(-60, 8),
    to_signed(-32, 8),
    to_signed(-6, 8),
    to_signed(7, 8),
    to_signed(4, 8),
    to_signed(-14, 8),
    to_signed(-38, 8),
    to_signed(-58, 8),
    to_signed(-70, 8),
    to_signed(-69, 8),
    to_signed(-57, 8),
    to_signed(-36, 8),
    to_signed(-11, 8),
    to_signed(14, 8),
    to_signed(35, 8),
    to_signed(46, 8),
    to_signed(48, 8),
    to_signed(41, 8),
    to_signed(32, 8),
    to_signed(22, 8),
    to_signed(14, 8),
    to_signed(6, 8),
    to_signed(0, 8),
    to_signed(-6, 8),
    to_signed(-15, 8),
    to_signed(-26, 8),
    to_signed(-36, 8),
    to_signed(-35, 8),
    to_signed(-22, 8),
    to_signed(-2, 8),
    to_signed(13, 8),
    to_signed(18, 8),
    to_signed(10, 8),
    to_signed(-8, 8),
    to_signed(-30, 8),
    to_signed(-47, 8),
    to_signed(-50, 8),
    to_signed(-40, 8),
    to_signed(-20, 8),
    to_signed(3, 8),
    to_signed(22, 8),
    to_signed(33, 8),
    to_signed(35, 8),
    to_signed(28, 8),
    to_signed(17, 8),
    to_signed(7, 8),
    to_signed(0, 8),
    to_signed(1, 8),
    to_signed(9, 8),
    to_signed(20, 8),
    to_signed(27, 8),
    to_signed(27, 8),
    to_signed(21, 8),
    to_signed(9, 8),
    to_signed(-5, 8),
    to_signed(-16, 8),
    to_signed(-19, 8),
    to_signed(-12, 8),
    to_signed(4, 8),
    to_signed(26, 8),
    to_signed(44, 8),
    to_signed(54, 8),
    to_signed(53, 8),
    to_signed(44, 8),
    to_signed(31, 8),
    to_signed(19, 8),
    to_signed(15, 8),
    to_signed(19, 8),
    to_signed(29, 8),
    to_signed(39, 8),
    to_signed(39, 8),
    to_signed(25, 8),
    to_signed(-2, 8),
    to_signed(-37, 8),
    to_signed(-67, 8),
    to_signed(-81, 8),
    to_signed(-77, 8),
    to_signed(-55, 8),
    to_signed(-25, 8),
    to_signed(1, 8),
    to_signed(12, 8),
    to_signed(7, 8),
    to_signed(-11, 8),
    to_signed(-33, 8),
    to_signed(-54, 8),
    to_signed(-65, 8),
    to_signed(-63, 8),
    to_signed(-47, 8),
    to_signed(-24, 8),
    to_signed(3, 8),
    to_signed(29, 8),
    to_signed(48, 8),
    to_signed(56, 8),
    to_signed(55, 8),
    to_signed(49, 8),
    to_signed(40, 8),
    to_signed(31, 8),
    to_signed(21, 8),
    to_signed(12, 8),
    to_signed(3, 8),
    to_signed(-8, 8),
    to_signed(-21, 8),
    to_signed(-34, 8),
    to_signed(-41, 8),
    to_signed(-39, 8),
    to_signed(-25, 8),
    to_signed(-5, 8),
    to_signed(12, 8),
    to_signed(18, 8),
    to_signed(9, 8),
    to_signed(-11, 8),
    to_signed(-35, 8),
    to_signed(-54, 8),
    to_signed(-62, 8),
    to_signed(-56, 8),
    to_signed(-42, 8),
    to_signed(-22, 8),
    to_signed(-3, 8),
    to_signed(9, 8),
    to_signed(14, 8),
    to_signed(13, 8),
    to_signed(11, 8),
    to_signed(6, 8),
    to_signed(3, 8),
    to_signed(3, 8),
    to_signed(9, 8),
    to_signed(16, 8),
    to_signed(20, 8),
    to_signed(21, 8),
    to_signed(19, 8),
    to_signed(13, 8),
    to_signed(5, 8),
    to_signed(-1, 8),
    to_signed(1, 8),
    to_signed(13, 8),
    to_signed(31, 8),
    to_signed(53, 8),
    to_signed(69, 8),
    to_signed(77, 8),
    to_signed(74, 8),
    to_signed(64, 8),
    to_signed(50, 8),
    to_signed(40, 8),
    to_signed(35, 8),
    to_signed(39, 8),
    to_signed(47, 8),
    to_signed(54, 8),
    to_signed(55, 8),
    to_signed(40, 8),
    to_signed(9, 8),
    to_signed(-31, 8),
    to_signed(-62, 8),
    to_signed(-75, 8),
    to_signed(-67, 8),
    to_signed(-43, 8),
    to_signed(-13, 8),
    to_signed(9, 8),
    to_signed(15, 8),
    to_signed(3, 8),
    to_signed(-21, 8),
    to_signed(-47, 8),
    to_signed(-70, 8),
    to_signed(-82, 8),
    to_signed(-79, 8),
    to_signed(-62, 8),
    to_signed(-38, 8),
    to_signed(-12, 8),
    to_signed(12, 8),
    to_signed(27, 8),
    to_signed(31, 8),
    to_signed(27, 8),
    to_signed(19, 8),
    to_signed(11, 8),
    to_signed(4, 8),
    to_signed(-4, 8),
    to_signed(-12, 8),
    to_signed(-22, 8),
    to_signed(-32, 8),
    to_signed(-42, 8),
    to_signed(-51, 8),
    to_signed(-55, 8),
    to_signed(-50, 8),
    to_signed(-33, 8),
    to_signed(-13, 8),
    to_signed(3, 8),
    to_signed(6, 8),
    to_signed(-1, 8),
    to_signed(-17, 8),
    to_signed(-36, 8),
    to_signed(-48, 8),
    to_signed(-47, 8),
    to_signed(-35, 8),
    to_signed(-15, 8),
    to_signed(6, 8),
    to_signed(22, 8),
    to_signed(33, 8),
    to_signed(38, 8),
    to_signed(39, 8),
    to_signed(38, 8),
    to_signed(35, 8),
    to_signed(32, 8),
    to_signed(32, 8),
    to_signed(33, 8),
    to_signed(33, 8),
    to_signed(32, 8),
    to_signed(31, 8),
    to_signed(28, 8),
    to_signed(21, 8),
    to_signed(11, 8),
    to_signed(5, 8),
    to_signed(7, 8),
    to_signed(18, 8),
    to_signed(35, 8),
    to_signed(51, 8),
    to_signed(60, 8),
    to_signed(60, 8),
    to_signed(51, 8),
    to_signed(38, 8),
    to_signed(23, 8),
    to_signed(11, 8),
    to_signed(8, 8),
    to_signed(14, 8),
    to_signed(24, 8),
    to_signed(33, 8),
    to_signed(32, 8),
    to_signed(14, 8),
    to_signed(-21, 8),
    to_signed(-65, 8),
    to_signed(-100, 8),
    to_signed(-115, 8),
    to_signed(-104, 8),
    to_signed(-75, 8),
    to_signed(-42, 8),
    to_signed(-19, 8),
    to_signed(-11, 8),
    to_signed(-16, 8),
    to_signed(-31, 8),
    to_signed(-50, 8),
    to_signed(-68, 8),
    to_signed(-77, 8),
    to_signed(-71, 8),
    to_signed(-55, 8),
    to_signed(-33, 8),
    to_signed(-11, 8),
    to_signed(10, 8),
    to_signed(25, 8),
    to_signed(32, 8),
    to_signed(33, 8),
    to_signed(33, 8),
    to_signed(33, 8),
    to_signed(31, 8),
    to_signed(25, 8),
    to_signed(16, 8),
    to_signed(3, 8),
    to_signed(-10, 8),
    to_signed(-22, 8),
    to_signed(-33, 8),
    to_signed(-38, 8),
    to_signed(-31, 8),
    to_signed(-15, 8),
    to_signed(7, 8),
    to_signed(23, 8),
    to_signed(28, 8),
    to_signed(20, 8),
    to_signed(3, 8),
    to_signed(-15, 8),
    to_signed(-27, 8),
    to_signed(-28, 8),
    to_signed(-21, 8),
    to_signed(-10, 8),
    to_signed(1, 8),
    to_signed(8, 8),
    to_signed(10, 8),
    to_signed(9, 8),
    to_signed(11, 8),
    to_signed(15, 8),
    to_signed(16, 8),
    to_signed(16, 8),
    to_signed(18, 8),
    to_signed(22, 8),
    to_signed(23, 8),
    to_signed(21, 8),
    to_signed(16, 8),
    to_signed(8, 8),
    to_signed(-2, 8),
    to_signed(-15, 8),
    to_signed(-24, 8),
    to_signed(-22, 8),
    to_signed(-6, 8),
    to_signed(18, 8),
    to_signed(41, 8),
    to_signed(56, 8),
    to_signed(62, 8),
    to_signed(59, 8),
    to_signed(48, 8),
    to_signed(33, 8),
    to_signed(21, 8),
    to_signed(15, 8),
    to_signed(18, 8),
    to_signed(26, 8),
    to_signed(33, 8),
    to_signed(30, 8),
    to_signed(10, 8),
    to_signed(-24, 8),
    to_signed(-62, 8),
    to_signed(-86, 8),
    to_signed(-86, 8),
    to_signed(-65, 8),
    to_signed(-33, 8),
    to_signed(-5, 8),
    to_signed(11, 8),
    to_signed(10, 8),
    to_signed(-6, 8),
    to_signed(-30, 8),
    to_signed(-54, 8),
    to_signed(-72, 8),
    to_signed(-75, 8),
    to_signed(-62, 8),
    to_signed(-37, 8),
    to_signed(-8, 8),
    to_signed(19, 8),
    to_signed(38, 8),
    to_signed(47, 8),
    to_signed(47, 8),
    to_signed(41, 8),
    to_signed(35, 8),
    to_signed(29, 8),
    to_signed(23, 8),
    to_signed(15, 8),
    to_signed(5, 8),
    to_signed(-7, 8),
    to_signed(-19, 8),
    to_signed(-31, 8),
    to_signed(-43, 8),
    to_signed(-50, 8),
    to_signed(-47, 8),
    to_signed(-32, 8),
    to_signed(-12, 8),
    to_signed(3, 8),
    to_signed(5, 8),
    to_signed(-5, 8),
    to_signed(-21, 8),
    to_signed(-36, 8),
    to_signed(-43, 8),
    to_signed(-41, 8),
    to_signed(-30, 8),
    to_signed(-14, 8),
    to_signed(3, 8),
    to_signed(17, 8),
    to_signed(25, 8),
    to_signed(31, 8),
    to_signed(35, 8),
    to_signed(36, 8),
    to_signed(34, 8),
    to_signed(29, 8),
    to_signed(26, 8),
    to_signed(25, 8),
    to_signed(23, 8),
    to_signed(20, 8),
    to_signed(14, 8),
    to_signed(4, 8),
    to_signed(-10, 8),
    to_signed(-23, 8),
    to_signed(-29, 8),
    to_signed(-23, 8),
    to_signed(-4, 8),
    to_signed(21, 8),
    to_signed(47, 8),
    to_signed(64, 8),
    to_signed(69, 8),
    to_signed(63, 8),
    to_signed(50, 8),
    to_signed(34, 8),
    to_signed(20, 8),
    to_signed(15, 8),
    to_signed(20, 8),
    to_signed(31, 8),
    to_signed(37, 8),
    to_signed(29, 8),
    to_signed(4, 8),
    to_signed(-32, 8),
    to_signed(-66, 8),
    to_signed(-82, 8),
    to_signed(-74, 8),
    to_signed(-46, 8),
    to_signed(-13, 8),
    to_signed(13, 8),
    to_signed(21, 8),
    to_signed(12, 8),
    to_signed(-9, 8),
    to_signed(-35, 8),
    to_signed(-60, 8),
    to_signed(-76, 8),
    to_signed(-73, 8),
    to_signed(-51, 8),
    to_signed(-18, 8),
    to_signed(12, 8),
    to_signed(36, 8),
    to_signed(49, 8),
    to_signed(52, 8),
    to_signed(45, 8),
    to_signed(35, 8),
    to_signed(25, 8),
    to_signed(16, 8),
    to_signed(8, 8),
    to_signed(0, 8),
    to_signed(-5, 8),
    to_signed(-9, 8),
    to_signed(-14, 8),
    to_signed(-21, 8),
    to_signed(-28, 8),
    to_signed(-29, 8),
    to_signed(-20, 8),
    to_signed(-2, 8),
    to_signed(15, 8),
    to_signed(25, 8),
    to_signed(21, 8),
    to_signed(6, 8),
    to_signed(-16, 8),
    to_signed(-36, 8),
    to_signed(-46, 8),
    to_signed(-44, 8),
    to_signed(-34, 8),
    to_signed(-21, 8),
    to_signed(-7, 8),
    to_signed(5, 8),
    to_signed(13, 8),
    to_signed(15, 8),
    to_signed(13, 8),
    to_signed(7, 8),
    to_signed(0, 8),
    to_signed(-6, 8),
    to_signed(-6, 8),
    to_signed(1, 8),
    to_signed(8, 8),
    to_signed(13, 8),
    to_signed(15, 8),
    to_signed(10, 8),
    to_signed(-1, 8),
    to_signed(-12, 8),
    to_signed(-17, 8),
    to_signed(-9, 8),
    to_signed(9, 8),
    to_signed(33, 8),
    to_signed(56, 8),
    to_signed(70, 8),
    to_signed(72, 8),
    to_signed(65, 8),
    to_signed(51, 8),
    to_signed(35, 8),
    to_signed(23, 8),
    to_signed(21, 8),
    to_signed(29, 8),
    to_signed(40, 8),
    to_signed(42, 8),
    to_signed(29, 8),
    to_signed(-1, 8),
    to_signed(-39, 8),
    to_signed(-70, 8),
    to_signed(-79, 8),
    to_signed(-66, 8),
    to_signed(-39, 8),
    to_signed(-9, 8),
    to_signed(13, 8),
    to_signed(21, 8),
    to_signed(12, 8),
    to_signed(-10, 8),
    to_signed(-36, 8),
    to_signed(-60, 8),
    to_signed(-72, 8),
    to_signed(-67, 8),
    to_signed(-45, 8),
    to_signed(-14, 8),
    to_signed(18, 8),
    to_signed(42, 8),
    to_signed(56, 8),
    to_signed(59, 8),
    to_signed(55, 8),
    to_signed(46, 8),
    to_signed(32, 8),
    to_signed(15, 8),
    to_signed(-3, 8),
    to_signed(-17, 8),
    to_signed(-25, 8),
    to_signed(-30, 8),
    to_signed(-34, 8),
    to_signed(-41, 8),
    to_signed(-47, 8),
    to_signed(-51, 8),
    to_signed(-45, 8),
    to_signed(-33, 8),
    to_signed(-20, 8),
    to_signed(-16, 8),
    to_signed(-21, 8),
    to_signed(-32, 8),
    to_signed(-43, 8),
    to_signed(-49, 8),
    to_signed(-47, 8),
    to_signed(-39, 8),
    to_signed(-27, 8),
    to_signed(-13, 8),
    to_signed(1, 8),
    to_signed(11, 8),
    to_signed(18, 8),
    to_signed(22, 8),
    to_signed(23, 8),
    to_signed(20, 8),
    to_signed(14, 8),
    to_signed(12, 8),
    to_signed(15, 8),
    to_signed(21, 8),
    to_signed(26, 8),
    to_signed(27, 8),
    to_signed(23, 8),
    to_signed(14, 8),
    to_signed(1, 8),
    to_signed(-8, 8),
    to_signed(-6, 8),
    to_signed(7, 8),
    to_signed(27, 8),
    to_signed(51, 8),
    to_signed(73, 8),
    to_signed(88, 8),
    to_signed(89, 8),
    to_signed(77, 8),
    to_signed(59, 8),
    to_signed(42, 8),
    to_signed(31, 8),
    to_signed(29, 8),
    to_signed(31, 8),
    to_signed(34, 8),
    to_signed(30, 8),
    to_signed(12, 8),
    to_signed(-21, 8),
    to_signed(-56, 8),
    to_signed(-78, 8),
    to_signed(-77, 8),
    to_signed(-58, 8),
    to_signed(-31, 8),
    to_signed(-6, 8),
    to_signed(9, 8),
    to_signed(10, 8),
    to_signed(-3, 8),
    to_signed(-27, 8),
    to_signed(-54, 8),
    to_signed(-77, 8),
    to_signed(-87, 8),
    to_signed(-79, 8),
    to_signed(-56, 8),
    to_signed(-28, 8),
    to_signed(-1, 8),
    to_signed(20, 8),
    to_signed(34, 8),
    to_signed(39, 8),
    to_signed(36, 8),
    to_signed(28, 8),
    to_signed(15, 8),
    to_signed(-2, 8),
    to_signed(-18, 8),
    to_signed(-28, 8),
    to_signed(-30, 8),
    to_signed(-28, 8),
    to_signed(-27, 8),
    to_signed(-29, 8),
    to_signed(-29, 8),
    to_signed(-23, 8),
    to_signed(-12, 8),
    to_signed(1, 8),
    to_signed(9, 8),
    to_signed(10, 8),
    to_signed(2, 8),
    to_signed(-13, 8),
    to_signed(-29, 8),
    to_signed(-39, 8),
    to_signed(-39, 8),
    to_signed(-33, 8),
    to_signed(-25, 8),
    to_signed(-16, 8),
    to_signed(-3, 8),
    to_signed(11, 8),
    to_signed(22, 8),
    to_signed(27, 8),
    to_signed(27, 8),
    to_signed(24, 8),
    to_signed(20, 8),
    to_signed(19, 8),
    to_signed(24, 8),
    to_signed(30, 8),
    to_signed(35, 8),
    to_signed(36, 8),
    to_signed(33, 8),
    to_signed(26, 8),
    to_signed(18, 8),
    to_signed(14, 8),
    to_signed(18, 8),
    to_signed(31, 8),
    to_signed(51, 8),
    to_signed(71, 8),
    to_signed(85, 8),
    to_signed(88, 8),
    to_signed(79, 8),
    to_signed(62, 8),
    to_signed(42, 8),
    to_signed(25, 8),
    to_signed(16, 8),
    to_signed(18, 8),
    to_signed(23, 8),
    to_signed(22, 8),
    to_signed(10, 8),
    to_signed(-16, 8),
    to_signed(-49, 8),
    to_signed(-79, 8),
    to_signed(-92, 8),
    to_signed(-84, 8),
    to_signed(-60, 8),
    to_signed(-30, 8),
    to_signed(-6, 8),
    to_signed(5, 8),
    to_signed(-1, 8),
    to_signed(-20, 8),
    to_signed(-46, 8),
    to_signed(-73, 8),
    to_signed(-90, 8),
    to_signed(-91, 8),
    to_signed(-74, 8),
    to_signed(-46, 8),
    to_signed(-16, 8),
    to_signed(12, 8),
    to_signed(33, 8),
    to_signed(44, 8),
    to_signed(43, 8),
    to_signed(36, 8),
    to_signed(27, 8),
    to_signed(16, 8),
    to_signed(2, 8),
    to_signed(-11, 8),
    to_signed(-19, 8),
    to_signed(-21, 8),
    to_signed(-21, 8),
    to_signed(-25, 8),
    to_signed(-30, 8),
    to_signed(-29, 8),
    to_signed(-20, 8),
    to_signed(-3, 8),
    to_signed(11, 8),
    to_signed(18, 8),
    to_signed(13, 8),
    to_signed(1, 8),
    to_signed(-15, 8),
    to_signed(-27, 8),
    to_signed(-31, 8),
    to_signed(-24, 8),
    to_signed(-11, 8),
    to_signed(7, 8),
    to_signed(26, 8),
    to_signed(42, 8),
    to_signed(53, 8),
    to_signed(57, 8),
    to_signed(54, 8),
    to_signed(44, 8),
    to_signed(33, 8),
    to_signed(25, 8),
    to_signed(24, 8),
    to_signed(29, 8),
    to_signed(33, 8),
    to_signed(32, 8),
    to_signed(24, 8),
    to_signed(11, 8),
    to_signed(-6, 8),
    to_signed(-22, 8),
    to_signed(-27, 8),
    to_signed(-20, 8),
    to_signed(-1, 8),
    to_signed(23, 8),
    to_signed(47, 8),
    to_signed(64, 8),
    to_signed(66, 8),
    to_signed(53, 8),
    to_signed(30, 8),
    to_signed(9, 8),
    to_signed(-3, 8),
    to_signed(-4, 8),
    to_signed(1, 8),
    to_signed(7, 8),
    to_signed(10, 8),
    to_signed(1, 8),
    to_signed(-23, 8),
    to_signed(-56, 8),
    to_signed(-82, 8),
    to_signed(-89, 8),
    to_signed(-77, 8),
    to_signed(-53, 8),
    to_signed(-25, 8),
    to_signed(-4, 8),
    to_signed(5, 8),
    to_signed(-2, 8),
    to_signed(-23, 8),
    to_signed(-49, 8),
    to_signed(-72, 8),
    to_signed(-83, 8),
    to_signed(-78, 8),
    to_signed(-55, 8),
    to_signed(-23, 8),
    to_signed(10, 8),
    to_signed(37, 8),
    to_signed(56, 8),
    to_signed(64, 8),
    to_signed(63, 8),
    to_signed(53, 8),
    to_signed(40, 8),
    to_signed(26, 8),
    to_signed(14, 8),
    to_signed(5, 8),
    to_signed(-1, 8),
    to_signed(-6, 8),
    to_signed(-11, 8),
    to_signed(-17, 8),
    to_signed(-21, 8),
    to_signed(-18, 8),
    to_signed(-7, 8),
    to_signed(7, 8),
    to_signed(17, 8),
    to_signed(17, 8),
    to_signed(6, 8),
    to_signed(-13, 8),
    to_signed(-34, 8),
    to_signed(-51, 8),
    to_signed(-58, 8),
    to_signed(-54, 8),
    to_signed(-42, 8),
    to_signed(-24, 8),
    to_signed(-7, 8),
    to_signed(7, 8),
    to_signed(15, 8),
    to_signed(15, 8),
    to_signed(8, 8),
    to_signed(-3, 8),
    to_signed(-13, 8),
    to_signed(-17, 8),
    to_signed(-14, 8),
    to_signed(-7, 8),
    to_signed(0, 8),
    to_signed(3, 8),
    to_signed(0, 8),
    to_signed(-6, 8),
    to_signed(-16, 8),
    to_signed(-22, 8),
    to_signed(-19, 8),
    to_signed(-6, 8),
    to_signed(16, 8),
    to_signed(40, 8),
    to_signed(61, 8),
    to_signed(70, 8),
    to_signed(67, 8),
    to_signed(53, 8),
    to_signed(34, 8),
    to_signed(19, 8),
    to_signed(12, 8),
    to_signed(15, 8),
    to_signed(24, 8),
    to_signed(32, 8),
    to_signed(30, 8),
    to_signed(14, 8),
    to_signed(-14, 8),
    to_signed(-44, 8),
    to_signed(-64, 8),
    to_signed(-67, 8),
    to_signed(-54, 8),
    to_signed(-30, 8),
    to_signed(-5, 8),
    to_signed(13, 8),
    to_signed(18, 8),
    to_signed(9, 8),
    to_signed(-14, 8),
    to_signed(-40, 8),
    to_signed(-62, 8),
    to_signed(-73, 8),
    to_signed(-67, 8),
    to_signed(-49, 8),
    to_signed(-21, 8),
    to_signed(8, 8),
    to_signed(35, 8),
    to_signed(55, 8),
    to_signed(62, 8),
    to_signed(59, 8),
    to_signed(49, 8),
    to_signed(35, 8),
    to_signed(18, 8),
    to_signed(0, 8),
    to_signed(-13, 8),
    to_signed(-21, 8),
    to_signed(-29, 8),
    to_signed(-39, 8),
    to_signed(-49, 8),
    to_signed(-52, 8),
    to_signed(-46, 8),
    to_signed(-35, 8),
    to_signed(-23, 8),
    to_signed(-17, 8),
    to_signed(-18, 8),
    to_signed(-25, 8),
    to_signed(-37, 8),
    to_signed(-50, 8),
    to_signed(-56, 8),
    to_signed(-54, 8),
    to_signed(-43, 8),
    to_signed(-26, 8),
    to_signed(-7, 8),
    to_signed(13, 8),
    to_signed(29, 8),
    to_signed(37, 8),
    to_signed(39, 8),
    to_signed(37, 8),
    to_signed(34, 8),
    to_signed(31, 8),
    to_signed(28, 8),
    to_signed(28, 8),
    to_signed(30, 8),
    to_signed(28, 8),
    to_signed(22, 8),
    to_signed(11, 8),
    to_signed(-3, 8),
    to_signed(-15, 8),
    to_signed(-18, 8),
    to_signed(-10, 8),
    to_signed(9, 8),
    to_signed(35, 8),
    to_signed(62, 8),
    to_signed(83, 8),
    to_signed(91, 8),
    to_signed(85, 8),
    to_signed(67, 8),
    to_signed(45, 8),
    to_signed(29, 8),
    to_signed(21, 8),
    to_signed(18, 8),
    to_signed(18, 8),
    to_signed(16, 8),
    to_signed(9, 8),
    to_signed(-10, 8),
    to_signed(-35, 8),
    to_signed(-58, 8),
    to_signed(-68, 8),
    to_signed(-62, 8),
    to_signed(-45, 8),
    to_signed(-27, 8),
    to_signed(-14, 8),
    to_signed(-10, 8),
    to_signed(-16, 8),
    to_signed(-33, 8),
    to_signed(-55, 8),
    to_signed(-74, 8),
    to_signed(-84, 8),
    to_signed(-79, 8),
    to_signed(-61, 8),
    to_signed(-33, 8),
    to_signed(-1, 8),
    to_signed(27, 8),
    to_signed(48, 8),
    to_signed(59, 8),
    to_signed(58, 8),
    to_signed(50, 8),
    to_signed(37, 8),
    to_signed(22, 8),
    to_signed(6, 8),
    to_signed(-6, 8),
    to_signed(-12, 8),
    to_signed(-15, 8),
    to_signed(-18, 8),
    to_signed(-22, 8),
    to_signed(-25, 8),
    to_signed(-23, 8),
    to_signed(-14, 8),
    to_signed(-3, 8),
    to_signed(4, 8),
    to_signed(4, 8),
    to_signed(-3, 8),
    to_signed(-15, 8),
    to_signed(-28, 8),
    to_signed(-38, 8),
    to_signed(-41, 8),
    to_signed(-38, 8),
    to_signed(-26, 8),
    to_signed(-9, 8),
    to_signed(8, 8),
    to_signed(23, 8),
    to_signed(33, 8),
    to_signed(37, 8),
    to_signed(35, 8),
    to_signed(29, 8),
    to_signed(24, 8),
    to_signed(21, 8),
    to_signed(21, 8),
    to_signed(25, 8),
    to_signed(28, 8),
    to_signed(28, 8),
    to_signed(25, 8),
    to_signed(19, 8),
    to_signed(9, 8),
    to_signed(0, 8),
    to_signed(0, 8),
    to_signed(10, 8),
    to_signed(26, 8),
    to_signed(45, 8),
    to_signed(63, 8),
    to_signed(72, 8),
    to_signed(71, 8),
    to_signed(60, 8),
    to_signed(45, 8),
    to_signed(30, 8),
    to_signed(21, 8),
    to_signed(19, 8),
    to_signed(19, 8),
    to_signed(18, 8),
    to_signed(13, 8),
    to_signed(-2, 8),
    to_signed(-26, 8),
    to_signed(-52, 8),
    to_signed(-66, 8),
    to_signed(-64, 8),
    to_signed(-46, 8),
    to_signed(-21, 8),
    to_signed(0, 8),
    to_signed(12, 8),
    to_signed(12, 8),
    to_signed(-1, 8),
    to_signed(-23, 8),
    to_signed(-48, 8),
    to_signed(-65, 8),
    to_signed(-68, 8),
    to_signed(-56, 8),
    to_signed(-31, 8),
    to_signed(0, 8),
    to_signed(30, 8),
    to_signed(53, 8),
    to_signed(68, 8),
    to_signed(71, 8),
    to_signed(65, 8),
    to_signed(55, 8),
    to_signed(42, 8),
    to_signed(26, 8),
    to_signed(9, 8),
    to_signed(-6, 8),
    to_signed(-16, 8),
    to_signed(-21, 8),
    to_signed(-26, 8),
    to_signed(-33, 8),
    to_signed(-39, 8),
    to_signed(-38, 8),
    to_signed(-29, 8),
    to_signed(-19, 8),
    to_signed(-14, 8),
    to_signed(-17, 8),
    to_signed(-26, 8),
    to_signed(-38, 8),
    to_signed(-51, 8),
    to_signed(-58, 8),
    to_signed(-59, 8),
    to_signed(-51, 8),
    to_signed(-34, 8),
    to_signed(-15, 8),
    to_signed(2, 8),
    to_signed(17, 8),
    to_signed(26, 8),
    to_signed(26, 8),
    to_signed(22, 8),
    to_signed(18, 8),
    to_signed(15, 8),
    to_signed(16, 8),
    to_signed(18, 8),
    to_signed(20, 8),
    to_signed(19, 8),
    to_signed(15, 8),
    to_signed(8, 8),
    to_signed(-1, 8),
    to_signed(-12, 8),
    to_signed(-16, 8),
    to_signed(-10, 8),
    to_signed(6, 8),
    to_signed(27, 8),
    to_signed(50, 8),
    to_signed(69, 8),
    to_signed(79, 8),
    to_signed(77, 8),
    to_signed(65, 8),
    to_signed(49, 8),
    to_signed(36, 8),
    to_signed(32, 8),
    to_signed(34, 8),
    to_signed(37, 8),
    to_signed(36, 8),
    to_signed(26, 8),
    to_signed(3, 8),
    to_signed(-27, 8),
    to_signed(-55, 8),
    to_signed(-70, 8),
    to_signed(-67, 8),
    to_signed(-50, 8),
    to_signed(-29, 8),
    to_signed(-13, 8),
    to_signed(-9, 8),
    to_signed(-15, 8),
    to_signed(-32, 8),
    to_signed(-55, 8),
    to_signed(-76, 8),
    to_signed(-89, 8),
    to_signed(-87, 8),
    to_signed(-70, 8),
    to_signed(-43, 8),
    to_signed(-13, 8),
    to_signed(13, 8),
    to_signed(31, 8),
    to_signed(40, 8),
    to_signed(40, 8),
    to_signed(34, 8),
    to_signed(26, 8),
    to_signed(15, 8),
    to_signed(2, 8),
    to_signed(-11, 8),
    to_signed(-21, 8),
    to_signed(-29, 8),
    to_signed(-35, 8),
    to_signed(-39, 8),
    to_signed(-44, 8),
    to_signed(-44, 8),
    to_signed(-37, 8),
    to_signed(-25, 8),
    to_signed(-13, 8),
    to_signed(-8, 8),
    to_signed(-12, 8),
    to_signed(-23, 8),
    to_signed(-35, 8),
    to_signed(-42, 8),
    to_signed(-43, 8),
    to_signed(-36, 8),
    to_signed(-21, 8),
    to_signed(0, 8),
    to_signed(20, 8),
    to_signed(36, 8),
    to_signed(46, 8),
    to_signed(47, 8),
    to_signed(43, 8),
    to_signed(36, 8),
    to_signed(29, 8),
    to_signed(25, 8),
    to_signed(27, 8),
    to_signed(33, 8),
    to_signed(40, 8),
    to_signed(40, 8),
    to_signed(33, 8),
    to_signed(20, 8),
    to_signed(5, 8),
    to_signed(-9, 8),
    to_signed(-17, 8),
    to_signed(-14, 8),
    to_signed(-2, 8),
    to_signed(20, 8),
    to_signed(43, 8),
    to_signed(61, 8),
    to_signed(68, 8),
    to_signed(61, 8),
    to_signed(46, 8),
    to_signed(29, 8),
    to_signed(15, 8),
    to_signed(9, 8),
    to_signed(8, 8),
    to_signed(10, 8),
    to_signed(8, 8),
    to_signed(-4, 8),
    to_signed(-27, 8),
    to_signed(-55, 8),
    to_signed(-76, 8),
    to_signed(-82, 8),
    to_signed(-70, 8),
    to_signed(-48, 8),
    to_signed(-25, 8),
    to_signed(-9, 8),
    to_signed(-4, 8),
    to_signed(-13, 8),
    to_signed(-35, 8),
    to_signed(-62, 8),
    to_signed(-83, 8),
    to_signed(-90, 8),
    to_signed(-77, 8),
    to_signed(-49, 8),
    to_signed(-13, 8),
    to_signed(23, 8),
    to_signed(53, 8),
    to_signed(71, 8),
    to_signed(76, 8),
    to_signed(72, 8),
    to_signed(65, 8),
    to_signed(54, 8),
    to_signed(42, 8),
    to_signed(28, 8),
    to_signed(17, 8),
    to_signed(9, 8),
    to_signed(4, 8),
    to_signed(-3, 8),
    to_signed(-11, 8),
    to_signed(-20, 8),
    to_signed(-24, 8),
    to_signed(-20, 8),
    to_signed(-14, 8),
    to_signed(-8, 8),
    to_signed(-7, 8),
    to_signed(-12, 8),
    to_signed(-22, 8),
    to_signed(-34, 8),
    to_signed(-45, 8),
    to_signed(-50, 8),
    to_signed(-46, 8),
    to_signed(-33, 8),
    to_signed(-15, 8),
    to_signed(4, 8),
    to_signed(21, 8),
    to_signed(31, 8),
    to_signed(31, 8),
    to_signed(27, 8),
    to_signed(20, 8),
    to_signed(13, 8),
    to_signed(8, 8),
    to_signed(4, 8),
    to_signed(3, 8),
    to_signed(2, 8),
    to_signed(1, 8),
    to_signed(-4, 8),
    to_signed(-13, 8),
    to_signed(-22, 8),
    to_signed(-28, 8),
    to_signed(-26, 8),
    to_signed(-18, 8),
    to_signed(-2, 8),
    to_signed(18, 8),
    to_signed(40, 8),
    to_signed(57, 8),
    to_signed(64, 8),
    to_signed(60, 8),
    to_signed(47, 8),
    to_signed(33, 8),
    to_signed(23, 8),
    to_signed(21, 8),
    to_signed(27, 8),
    to_signed(32, 8),
    to_signed(29, 8),
    to_signed(12, 8),
    to_signed(-14, 8),
    to_signed(-40, 8),
    to_signed(-55, 8),
    to_signed(-52, 8),
    to_signed(-35, 8),
    to_signed(-13, 8),
    to_signed(7, 8),
    to_signed(19, 8),
    to_signed(17, 8),
    to_signed(0, 8),
    to_signed(-25, 8),
    to_signed(-49, 8),
    to_signed(-65, 8),
    to_signed(-68, 8),
    to_signed(-54, 8),
    to_signed(-28, 8),
    to_signed(4, 8),
    to_signed(33, 8),
    to_signed(54, 8),
    to_signed(62, 8),
    to_signed(59, 8),
    to_signed(51, 8),
    to_signed(38, 8),
    to_signed(23, 8),
    to_signed(7, 8),
    to_signed(-7, 8),
    to_signed(-16, 8),
    to_signed(-22, 8),
    to_signed(-25, 8),
    to_signed(-30, 8),
    to_signed(-37, 8),
    to_signed(-40, 8),
    to_signed(-37, 8),
    to_signed(-28, 8),
    to_signed(-18, 8),
    to_signed(-14, 8),
    to_signed(-18, 8),
    to_signed(-28, 8),
    to_signed(-42, 8),
    to_signed(-54, 8),
    to_signed(-62, 8),
    to_signed(-61, 8),
    to_signed(-50, 8),
    to_signed(-32, 8),
    to_signed(-13, 8),
    to_signed(6, 8),
    to_signed(18, 8),
    to_signed(22, 8),
    to_signed(18, 8),
    to_signed(12, 8),
    to_signed(7, 8),
    to_signed(5, 8),
    to_signed(7, 8),
    to_signed(12, 8),
    to_signed(18, 8),
    to_signed(25, 8),
    to_signed(28, 8),
    to_signed(25, 8),
    to_signed(14, 8),
    to_signed(2, 8),
    to_signed(-6, 8),
    to_signed(-6, 8),
    to_signed(4, 8),
    to_signed(20, 8),
    to_signed(38, 8),
    to_signed(56, 8),
    to_signed(69, 8),
    to_signed(71, 8),
    to_signed(62, 8),
    to_signed(47, 8),
    to_signed(32, 8),
    to_signed(24, 8),
    to_signed(24, 8),
    to_signed(29, 8),
    to_signed(33, 8),
    to_signed(27, 8),
    to_signed(8, 8),
    to_signed(-21, 8),
    to_signed(-49, 8),
    to_signed(-64, 8),
    to_signed(-59, 8),
    to_signed(-41, 8),
    to_signed(-20, 8),
    to_signed(-3, 8),
    to_signed(7, 8),
    to_signed(4, 8),
    to_signed(-12, 8),
    to_signed(-35, 8),
    to_signed(-58, 8),
    to_signed(-73, 8),
    to_signed(-71, 8),
    to_signed(-52, 8),
    to_signed(-25, 8),
    to_signed(3, 8),
    to_signed(28, 8),
    to_signed(44, 8),
    to_signed(49, 8),
    to_signed(48, 8),
    to_signed(43, 8),
    to_signed(35, 8),
    to_signed(24, 8),
    to_signed(11, 8),
    to_signed(-3, 8),
    to_signed(-14, 8),
    to_signed(-21, 8),
    to_signed(-25, 8),
    to_signed(-29, 8),
    to_signed(-31, 8),
    to_signed(-29, 8),
    to_signed(-22, 8),
    to_signed(-10, 8),
    to_signed(1, 8),
    to_signed(5, 8),
    to_signed(-3, 8),
    to_signed(-18, 8),
    to_signed(-34, 8),
    to_signed(-48, 8),
    to_signed(-54, 8),
    to_signed(-49, 8),
    to_signed(-34, 8),
    to_signed(-14, 8),
    to_signed(8, 8),
    to_signed(27, 8),
    to_signed(37, 8),
    to_signed(34, 8),
    to_signed(26, 8),
    to_signed(16, 8),
    to_signed(10, 8),
    to_signed(9, 8),
    to_signed(13, 8),
    to_signed(18, 8),
    to_signed(23, 8),
    to_signed(27, 8),
    to_signed(27, 8),
    to_signed(22, 8),
    to_signed(13, 8),
    to_signed(3, 8),
    to_signed(-3, 8),
    to_signed(0, 8),
    to_signed(12, 8),
    to_signed(30, 8),
    to_signed(47, 8),
    to_signed(61, 8),
    to_signed(67, 8),
    to_signed(65, 8),
    to_signed(54, 8),
    to_signed(41, 8),
    to_signed(29, 8),
    to_signed(25, 8),
    to_signed(31, 8),
    to_signed(42, 8),
    to_signed(46, 8),
    to_signed(36, 8),
    to_signed(10, 8),
    to_signed(-25, 8),
    to_signed(-56, 8),
    to_signed(-69, 8),
    to_signed(-62, 8),
    to_signed(-43, 8),
    to_signed(-20, 8),
    to_signed(1, 8),
    to_signed(13, 8),
    to_signed(10, 8),
    to_signed(-6, 8),
    to_signed(-29, 8),
    to_signed(-52, 8),
    to_signed(-66, 8),
    to_signed(-64, 8),
    to_signed(-47, 8),
    to_signed(-20, 8),
    to_signed(9, 8),
    to_signed(35, 8),
    to_signed(51, 8),
    to_signed(57, 8),
    to_signed(57, 8),
    to_signed(54, 8),
    to_signed(47, 8),
    to_signed(37, 8),
    to_signed(25, 8),
    to_signed(12, 8),
    to_signed(0, 8),
    to_signed(-10, 8),
    to_signed(-21, 8),
    to_signed(-34, 8),
    to_signed(-44, 8),
    to_signed(-46, 8),
    to_signed(-38, 8),
    to_signed(-24, 8),
    to_signed(-11, 8),
    to_signed(-6, 8),
    to_signed(-10, 8),
    to_signed(-21, 8),
    to_signed(-35, 8),
    to_signed(-47, 8),
    to_signed(-52, 8),
    to_signed(-45, 8),
    to_signed(-31, 8),
    to_signed(-14, 8),
    to_signed(4, 8),
    to_signed(18, 8),
    to_signed(26, 8),
    to_signed(28, 8),
    to_signed(26, 8),
    to_signed(22, 8),
    to_signed(19, 8),
    to_signed(20, 8),
    to_signed(23, 8),
    to_signed(26, 8),
    to_signed(27, 8),
    to_signed(25, 8),
    to_signed(19, 8),
    to_signed(9, 8),
    to_signed(0, 8),
    to_signed(-8, 8),
    to_signed(-12, 8),
    to_signed(-6, 8),
    to_signed(11, 8),
    to_signed(35, 8),
    to_signed(56, 8),
    to_signed(70, 8),
    to_signed(73, 8),
    to_signed(66, 8),
    to_signed(53, 8),
    to_signed(38, 8),
    to_signed(24, 8),
    to_signed(19, 8),
    to_signed(23, 8),
    to_signed(31, 8),
    to_signed(34, 8),
    to_signed(25, 8),
    to_signed(1, 8),
    to_signed(-30, 8),
    to_signed(-56, 8),
    to_signed(-65, 8),
    to_signed(-57, 8),
    to_signed(-40, 8),
    to_signed(-20, 8),
    to_signed(-3, 8),
    to_signed(2, 8),
    to_signed(-8, 8),
    to_signed(-30, 8),
    to_signed(-55, 8),
    to_signed(-78, 8),
    to_signed(-88, 8),
    to_signed(-80, 8),
    to_signed(-58, 8),
    to_signed(-28, 8),
    to_signed(1, 8),
    to_signed(22, 8),
    to_signed(32, 8),
    to_signed(33, 8),
    to_signed(29, 8),
    to_signed(24, 8),
    to_signed(18, 8),
    to_signed(11, 8),
    to_signed(3, 8),
    to_signed(-5, 8),
    to_signed(-11, 8),
    to_signed(-18, 8),
    to_signed(-25, 8),
    to_signed(-33, 8),
    to_signed(-37, 8),
    to_signed(-35, 8),
    to_signed(-24, 8),
    to_signed(-10, 8),
    to_signed(1, 8),
    to_signed(3, 8),
    to_signed(-3, 8),
    to_signed(-16, 8),
    to_signed(-33, 8),
    to_signed(-47, 8),
    to_signed(-50, 8),
    to_signed(-41, 8),
    to_signed(-24, 8),
    to_signed(-4, 8),
    to_signed(15, 8),
    to_signed(30, 8),
    to_signed(38, 8),
    to_signed(38, 8),
    to_signed(33, 8),
    to_signed(25, 8),
    to_signed(17, 8),
    to_signed(14, 8),
    to_signed(15, 8),
    to_signed(17, 8),
    to_signed(18, 8),
    to_signed(15, 8),
    to_signed(8, 8),
    to_signed(-4, 8),
    to_signed(-16, 8),
    to_signed(-25, 8),
    to_signed(-26, 8),
    to_signed(-18, 8),
    to_signed(0, 8),
    to_signed(22, 8),
    to_signed(41, 8),
    to_signed(51, 8),
    to_signed(48, 8),
    to_signed(37, 8),
    to_signed(21, 8),
    to_signed(6, 8),
    to_signed(-3, 8),
    to_signed(-1, 8),
    to_signed(9, 8),
    to_signed(20, 8),
    to_signed(24, 8),
    to_signed(14, 8),
    to_signed(-10, 8),
    to_signed(-43, 8),
    to_signed(-68, 8),
    to_signed(-75, 8),
    to_signed(-66, 8),
    to_signed(-47, 8),
    to_signed(-25, 8),
    to_signed(-6, 8),
    to_signed(0, 8),
    to_signed(-7, 8),
    to_signed(-25, 8),
    to_signed(-46, 8),
    to_signed(-64, 8),
    to_signed(-68, 8),
    to_signed(-57, 8),
    to_signed(-34, 8),
    to_signed(-5, 8),
    to_signed(23, 8),
    to_signed(42, 8),
    to_signed(51, 8),
    to_signed(51, 8),
    to_signed(46, 8),
    to_signed(39, 8),
    to_signed(31, 8),
    to_signed(22, 8),
    to_signed(14, 8),
    to_signed(6, 8),
    to_signed(-1, 8),
    to_signed(-10, 8),
    to_signed(-20, 8),
    to_signed(-31, 8),
    to_signed(-39, 8),
    to_signed(-38, 8),
    to_signed(-29, 8),
    to_signed(-15, 8),
    to_signed(-5, 8),
    to_signed(-6, 8),
    to_signed(-14, 8),
    to_signed(-27, 8),
    to_signed(-41, 8),
    to_signed(-52, 8),
    to_signed(-54, 8),
    to_signed(-45, 8),
    to_signed(-29, 8),
    to_signed(-11, 8),
    to_signed(5, 8),
    to_signed(14, 8),
    to_signed(15, 8),
    to_signed(12, 8),
    to_signed(8, 8),
    to_signed(3, 8),
    to_signed(-2, 8),
    to_signed(-3, 8),
    to_signed(2, 8),
    to_signed(9, 8),
    to_signed(15, 8),
    to_signed(14, 8),
    to_signed(4, 8),
    to_signed(-10, 8),
    to_signed(-22, 8),
    to_signed(-26, 8),
    to_signed(-21, 8),
    to_signed(-6, 8),
    to_signed(16, 8),
    to_signed(41, 8),
    to_signed(62, 8),
    to_signed(72, 8),
    to_signed(67, 8),
    to_signed(53, 8),
    to_signed(38, 8),
    to_signed(27, 8),
    to_signed(26, 8),
    to_signed(35, 8),
    to_signed(49, 8),
    to_signed(59, 8),
    to_signed(58, 8),
    to_signed(43, 8),
    to_signed(12, 8),
    to_signed(-25, 8),
    to_signed(-51, 8),
    to_signed(-57, 8),
    to_signed(-46, 8),
    to_signed(-27, 8),
    to_signed(-7, 8),
    to_signed(6, 8),
    to_signed(7, 8),
    to_signed(-6, 8),
    to_signed(-28, 8),
    to_signed(-52, 8),
    to_signed(-69, 8),
    to_signed(-72, 8),
    to_signed(-60, 8),
    to_signed(-40, 8),
    to_signed(-19, 8),
    to_signed(-1, 8),
    to_signed(12, 8),
    to_signed(19, 8),
    to_signed(21, 8),
    to_signed(21, 8),
    to_signed(19, 8),
    to_signed(17, 8),
    to_signed(12, 8),
    to_signed(3, 8),
    to_signed(-8, 8),
    to_signed(-20, 8),
    to_signed(-31, 8),
    to_signed(-43, 8),
    to_signed(-53, 8),
    to_signed(-57, 8),
    to_signed(-52, 8),
    to_signed(-38, 8),
    to_signed(-20, 8),
    to_signed(-9, 8),
    to_signed(-8, 8),
    to_signed(-17, 8),
    to_signed(-28, 8),
    to_signed(-38, 8),
    to_signed(-44, 8),
    to_signed(-42, 8),
    to_signed(-31, 8),
    to_signed(-13, 8),
    to_signed(8, 8),
    to_signed(26, 8),
    to_signed(35, 8),
    to_signed(35, 8),
    to_signed(32, 8),
    to_signed(29, 8),
    to_signed(26, 8),
    to_signed(24, 8),
    to_signed(28, 8),
    to_signed(37, 8),
    to_signed(47, 8),
    to_signed(50, 8),
    to_signed(42, 8),
    to_signed(26, 8),
    to_signed(7, 8),
    to_signed(-7, 8),
    to_signed(-11, 8),
    to_signed(-5, 8),
    to_signed(11, 8),
    to_signed(33, 8),
    to_signed(56, 8),
    to_signed(72, 8),
    to_signed(75, 8),
    to_signed(64, 8),
    to_signed(46, 8),
    to_signed(28, 8),
    to_signed(16, 8),
    to_signed(13, 8),
    to_signed(18, 8),
    to_signed(26, 8),
    to_signed(26, 8),
    to_signed(13, 8),
    to_signed(-12, 8),
    to_signed(-46, 8),
    to_signed(-74, 8),
    to_signed(-85, 8),
    to_signed(-77, 8),
    to_signed(-57, 8),
    to_signed(-34, 8),
    to_signed(-17, 8),
    to_signed(-13, 8),
    to_signed(-25, 8),
    to_signed(-48, 8),
    to_signed(-71, 8),
    to_signed(-89, 8),
    to_signed(-93, 8),
    to_signed(-83, 8),
    to_signed(-60, 8),
    to_signed(-32, 8),
    to_signed(-6, 8),
    to_signed(15, 8),
    to_signed(27, 8),
    to_signed(31, 8),
    to_signed(31, 8),
    to_signed(27, 8),
    to_signed(22, 8),
    to_signed(18, 8),
    to_signed(13, 8),
    to_signed(7, 8),
    to_signed(1, 8),
    to_signed(-3, 8),
    to_signed(-8, 8),
    to_signed(-14, 8),
    to_signed(-19, 8),
    to_signed(-17, 8),
    to_signed(-6, 8),
    to_signed(13, 8),
    to_signed(29, 8),
    to_signed(34, 8),
    to_signed(27, 8),
    to_signed(10, 8),
    to_signed(-6, 8),
    to_signed(-18, 8),
    to_signed(-21, 8),
    to_signed(-16, 8),
    to_signed(-4, 8),
    to_signed(11, 8),
    to_signed(27, 8),
    to_signed(38, 8),
    to_signed(40, 8),
    to_signed(34, 8),
    to_signed(25, 8),
    to_signed(15, 8),
    to_signed(7, 8),
    to_signed(4, 8),
    to_signed(7, 8),
    to_signed(14, 8),
    to_signed(20, 8),
    to_signed(19, 8),
    to_signed(12, 8),
    to_signed(0, 8),
    to_signed(-11, 8),
    to_signed(-18, 8),
    to_signed(-15, 8),
    to_signed(-4, 8),
    to_signed(13, 8),
    to_signed(31, 8),
    to_signed(44, 8),
    to_signed(49, 8),
    to_signed(44, 8),
    to_signed(30, 8),
    to_signed(15, 8),
    to_signed(2, 8),
    to_signed(-4, 8),
    to_signed(-1, 8),
    to_signed(9, 8),
    to_signed(14, 8),
    to_signed(6, 8),
    to_signed(-16, 8),
    to_signed(-47, 8),
    to_signed(-79, 8),
    to_signed(-97, 8),
    to_signed(-95, 8),
    to_signed(-75, 8),
    to_signed(-46, 8),
    to_signed(-17, 8),
    to_signed(0, 8),
    to_signed(0, 8),
    to_signed(-16, 8),
    to_signed(-39, 8),
    to_signed(-58, 8),
    to_signed(-67, 8),
    to_signed(-61, 8),
    to_signed(-41, 8),
    to_signed(-11, 8),
    to_signed(21, 8),
    to_signed(45, 8),
    to_signed(60, 8),
    to_signed(65, 8),
    to_signed(64, 8),
    to_signed(60, 8),
    to_signed(53, 8),
    to_signed(44, 8),
    to_signed(36, 8),
    to_signed(28, 8),
    to_signed(20, 8),
    to_signed(12, 8),
    to_signed(5, 8),
    to_signed(-3, 8),
    to_signed(-11, 8),
    to_signed(-17, 8),
    to_signed(-18, 8),
    to_signed(-11, 8),
    to_signed(-1, 8),
    to_signed(6, 8),
    to_signed(5, 8),
    to_signed(-7, 8),
    to_signed(-23, 8),
    to_signed(-36, 8),
    to_signed(-41, 8),
    to_signed(-36, 8),
    to_signed(-25, 8),
    to_signed(-11, 8),
    to_signed(4, 8),
    to_signed(20, 8),
    to_signed(31, 8),
    to_signed(33, 8),
    to_signed(26, 8),
    to_signed(16, 8),
    to_signed(8, 8),
    to_signed(3, 8),
    to_signed(2, 8),
    to_signed(4, 8),
    to_signed(7, 8),
    to_signed(7, 8),
    to_signed(1, 8),
    to_signed(-11, 8),
    to_signed(-23, 8),
    to_signed(-33, 8),
    to_signed(-36, 8),
    to_signed(-27, 8),
    to_signed(-11, 8),
    to_signed(9, 8),
    to_signed(27, 8),
    to_signed(39, 8),
    to_signed(42, 8),
    to_signed(35, 8),
    to_signed(23, 8),
    to_signed(11, 8),
    to_signed(4, 8),
    to_signed(6, 8),
    to_signed(17, 8),
    to_signed(31, 8),
    to_signed(40, 8),
    to_signed(35, 8),
    to_signed(15, 8),
    to_signed(-13, 8),
    to_signed(-38, 8),
    to_signed(-49, 8),
    to_signed(-42, 8),
    to_signed(-21, 8),
    to_signed(4, 8),
    to_signed(23, 8),
    to_signed(30, 8),
    to_signed(23, 8),
    to_signed(6, 8),
    to_signed(-14, 8),
    to_signed(-28, 8),
    to_signed(-33, 8),
    to_signed(-26, 8),
    to_signed(-9, 8),
    to_signed(10, 8),
    to_signed(27, 8),
    to_signed(38, 8),
    to_signed(43, 8),
    to_signed(42, 8),
    to_signed(40, 8),
    to_signed(36, 8),
    to_signed(30, 8),
    to_signed(22, 8),
    to_signed(14, 8),
    to_signed(7, 8),
    to_signed(1, 8),
    to_signed(-7, 8),
    to_signed(-15, 8),
    to_signed(-21, 8),
    to_signed(-24, 8),
    to_signed(-22, 8),
    to_signed(-14, 8),
    to_signed(-1, 8),
    to_signed(9, 8),
    to_signed(11, 8),
    to_signed(2, 8),
    to_signed(-17, 8),
    to_signed(-39, 8),
    to_signed(-56, 8),
    to_signed(-59, 8),
    to_signed(-51, 8),
    to_signed(-38, 8),
    to_signed(-24, 8),
    to_signed(-13, 8),
    to_signed(-5, 8),
    to_signed(-2, 8),
    to_signed(-6, 8),
    to_signed(-15, 8),
    to_signed(-23, 8),
    to_signed(-27, 8),
    to_signed(-24, 8),
    to_signed(-16, 8),
    to_signed(-5, 8),
    to_signed(5, 8),
    to_signed(13, 8),
    to_signed(15, 8),
    to_signed(12, 8),
    to_signed(7, 8),
    to_signed(4, 8),
    to_signed(7, 8),
    to_signed(18, 8),
    to_signed(35, 8),
    to_signed(56, 8),
    to_signed(74, 8),
    to_signed(84, 8),
    to_signed(84, 8),
    to_signed(75, 8),
    to_signed(61, 8),
    to_signed(49, 8),
    to_signed(45, 8),
    to_signed(50, 8),
    to_signed(59, 8),
    to_signed(67, 8),
    to_signed(67, 8),
    to_signed(52, 8),
    to_signed(22, 8),
    to_signed(-15, 8),
    to_signed(-45, 8),
    to_signed(-59, 8),
    to_signed(-54, 8),
    to_signed(-35, 8),
    to_signed(-10, 8),
    to_signed(11, 8),
    to_signed(20, 8),
    to_signed(15, 8),
    to_signed(-1, 8),
    to_signed(-23, 8),
    to_signed(-44, 8),
    to_signed(-55, 8),
    to_signed(-55, 8),
    to_signed(-45, 8),
    to_signed(-30, 8),
    to_signed(-16, 8),
    to_signed(-4, 8),
    to_signed(5, 8),
    to_signed(8, 8),
    to_signed(9, 8),
    to_signed(10, 8),
    to_signed(8, 8),
    to_signed(2, 8),
    to_signed(-7, 8),
    to_signed(-18, 8),
    to_signed(-30, 8),
    to_signed(-41, 8),
    to_signed(-51, 8),
    to_signed(-57, 8),
    to_signed(-59, 8),
    to_signed(-54, 8),
    to_signed(-41, 8),
    to_signed(-25, 8),
    to_signed(-12, 8),
    to_signed(-6, 8),
    to_signed(-8, 8),
    to_signed(-17, 8),
    to_signed(-30, 8),
    to_signed(-39, 8),
    to_signed(-40, 8),
    to_signed(-33, 8),
    to_signed(-21, 8),
    to_signed(-6, 8),
    to_signed(8, 8),
    to_signed(17, 8),
    to_signed(23, 8),
    to_signed(27, 8),
    to_signed(27, 8),
    to_signed(25, 8),
    to_signed(24, 8),
    to_signed(29, 8),
    to_signed(38, 8),
    to_signed(47, 8),
    to_signed(51, 8),
    to_signed(48, 8),
    to_signed(41, 8),
    to_signed(30, 8),
    to_signed(21, 8),
    to_signed(16, 8),
    to_signed(18, 8),
    to_signed(27, 8),
    to_signed(43, 8),
    to_signed(64, 8),
    to_signed(81, 8),
    to_signed(87, 8),
    to_signed(80, 8),
    to_signed(64, 8),
    to_signed(45, 8),
    to_signed(28, 8),
    to_signed(19, 8),
    to_signed(20, 8),
    to_signed(27, 8),
    to_signed(34, 8),
    to_signed(33, 8),
    to_signed(16, 8),
    to_signed(-16, 8),
    to_signed(-50, 8),
    to_signed(-73, 8),
    to_signed(-78, 8),
    to_signed(-68, 8),
    to_signed(-45, 8),
    to_signed(-19, 8),
    to_signed(0, 8),
    to_signed(2, 8),
    to_signed(-12, 8),
    to_signed(-37, 8),
    to_signed(-63, 8),
    to_signed(-82, 8),
    to_signed(-88, 8),
    to_signed(-80, 8),
    to_signed(-61, 8),
    to_signed(-37, 8),
    to_signed(-13, 8),
    to_signed(6, 8),
    to_signed(14, 8),
    to_signed(11, 8),
    to_signed(7, 8),
    to_signed(7, 8),
    to_signed(7, 8),
    to_signed(3, 8),
    to_signed(-2, 8),
    to_signed(-5, 8),
    to_signed(-6, 8),
    to_signed(-7, 8),
    to_signed(-9, 8),
    to_signed(-11, 8),
    to_signed(-9, 8),
    to_signed(0, 8),
    to_signed(15, 8),
    to_signed(29, 8),
    to_signed(37, 8),
    to_signed(39, 8),
    to_signed(33, 8),
    to_signed(19, 8),
    to_signed(0, 8),
    to_signed(-14, 8),
    to_signed(-18, 8),
    to_signed(-11, 8),
    to_signed(4, 8),
    to_signed(18, 8),
    to_signed(29, 8),
    to_signed(34, 8),
    to_signed(36, 8),
    to_signed(33, 8),
    to_signed(27, 8),
    to_signed(18, 8),
    to_signed(11, 8),
    to_signed(13, 8),
    to_signed(21, 8),
    to_signed(28, 8),
    to_signed(30, 8),
    to_signed(30, 8),
    to_signed(25, 8),
    to_signed(15, 8),
    to_signed(4, 8),
    to_signed(-2, 8),
    to_signed(-1, 8),
    to_signed(5, 8),
    to_signed(18, 8),
    to_signed(35, 8),
    to_signed(50, 8),
    to_signed(55, 8),
    to_signed(51, 8),
    to_signed(39, 8),
    to_signed(21, 8),
    to_signed(6, 8),
    to_signed(-1, 8),
    to_signed(3, 8),
    to_signed(12, 8),
    to_signed(19, 8),
    to_signed(17, 8),
    to_signed(0, 8),
    to_signed(-29, 8),
    to_signed(-62, 8),
    to_signed(-85, 8),
    to_signed(-90, 8),
    to_signed(-77, 8),
    to_signed(-52, 8),
    to_signed(-25, 8),
    to_signed(-7, 8),
    to_signed(-3, 8),
    to_signed(-15, 8),
    to_signed(-36, 8),
    to_signed(-58, 8),
    to_signed(-73, 8),
    to_signed(-75, 8),
    to_signed(-62, 8),
    to_signed(-38, 8),
    to_signed(-12, 8),
    to_signed(11, 8),
    to_signed(28, 8),
    to_signed(35, 8),
    to_signed(32, 8),
    to_signed(29, 8),
    to_signed(31, 8),
    to_signed(33, 8),
    to_signed(29, 8),
    to_signed(19, 8),
    to_signed(8, 8),
    to_signed(-2, 8),
    to_signed(-11, 8),
    to_signed(-17, 8),
    to_signed(-21, 8),
    to_signed(-21, 8),
    to_signed(-15, 8),
    to_signed(-2, 8),
    to_signed(10, 8),
    to_signed(15, 8),
    to_signed(12, 8),
    to_signed(2, 8),
    to_signed(-14, 8),
    to_signed(-31, 8),
    to_signed(-44, 8),
    to_signed(-47, 8),
    to_signed(-39, 8),
    to_signed(-24, 8),
    to_signed(-7, 8),
    to_signed(6, 8),
    to_signed(12, 8),
    to_signed(13, 8),
    to_signed(11, 8),
    to_signed(5, 8),
    to_signed(-4, 8),
    to_signed(-11, 8),
    to_signed(-10, 8),
    to_signed(-4, 8),
    to_signed(1, 8),
    to_signed(2, 8),
    to_signed(2, 8),
    to_signed(0, 8),
    to_signed(-6, 8),
    to_signed(-15, 8),
    to_signed(-18, 8),
    to_signed(-14, 8),
    to_signed(-5, 8),
    to_signed(11, 8),
    to_signed(30, 8),
    to_signed(45, 8),
    to_signed(51, 8),
    to_signed(48, 8),
    to_signed(38, 8),
    to_signed(22, 8),
    to_signed(7, 8),
    to_signed(2, 8),
    to_signed(10, 8),
    to_signed(26, 8),
    to_signed(40, 8),
    to_signed(45, 8),
    to_signed(33, 8),
    to_signed(3, 8),
    to_signed(-35, 8),
    to_signed(-67, 8),
    to_signed(-80, 8),
    to_signed(-71, 8),
    to_signed(-47, 8),
    to_signed(-20, 8),
    to_signed(1, 8),
    to_signed(8, 8),
    to_signed(-1, 8),
    to_signed(-21, 8),
    to_signed(-45, 8),
    to_signed(-66, 8),
    to_signed(-74, 8),
    to_signed(-66, 8),
    to_signed(-46, 8),
    to_signed(-24, 8),
    to_signed(-5, 8),
    to_signed(9, 8),
    to_signed(14, 8),
    to_signed(11, 8),
    to_signed(7, 8),
    to_signed(8, 8),
    to_signed(12, 8),
    to_signed(13, 8),
    to_signed(10, 8),
    to_signed(3, 8),
    to_signed(-8, 8),
    to_signed(-19, 8),
    to_signed(-28, 8),
    to_signed(-35, 8),
    to_signed(-37, 8),
    to_signed(-33, 8),
    to_signed(-19, 8),
    to_signed(-2, 8),
    to_signed(8, 8),
    to_signed(7, 8),
    to_signed(-3, 8),
    to_signed(-19, 8),
    to_signed(-36, 8),
    to_signed(-49, 8),
    to_signed(-52, 8),
    to_signed(-44, 8),
    to_signed(-29, 8),
    to_signed(-11, 8),
    to_signed(4, 8),
    to_signed(13, 8),
    to_signed(16, 8),
    to_signed(16, 8),
    to_signed(15, 8),
    to_signed(12, 8),
    to_signed(8, 8),
    to_signed(9, 8),
    to_signed(14, 8),
    to_signed(20, 8),
    to_signed(22, 8),
    to_signed(21, 8),
    to_signed(17, 8),
    to_signed(7, 8),
    to_signed(-5, 8),
    to_signed(-13, 8),
    to_signed(-12, 8),
    to_signed(-4, 8),
    to_signed(10, 8),
    to_signed(29, 8),
    to_signed(45, 8),
    to_signed(52, 8),
    to_signed(50, 8),
    to_signed(40, 8),
    to_signed(26, 8),
    to_signed(12, 8),
    to_signed(5, 8),
    to_signed(10, 8),
    to_signed(24, 8),
    to_signed(39, 8),
    to_signed(47, 8),
    to_signed(41, 8),
    to_signed(16, 8),
    to_signed(-21, 8),
    to_signed(-56, 8),
    to_signed(-73, 8),
    to_signed(-67, 8),
    to_signed(-44, 8),
    to_signed(-16, 8),
    to_signed(7, 8),
    to_signed(17, 8),
    to_signed(10, 8),
    to_signed(-11, 8),
    to_signed(-37, 8),
    to_signed(-60, 8),
    to_signed(-72, 8),
    to_signed(-68, 8),
    to_signed(-50, 8),
    to_signed(-26, 8),
    to_signed(-6, 8),
    to_signed(8, 8),
    to_signed(15, 8),
    to_signed(14, 8),
    to_signed(8, 8),
    to_signed(4, 8),
    to_signed(5, 8),
    to_signed(8, 8),
    to_signed(7, 8),
    to_signed(2, 8),
    to_signed(-7, 8),
    to_signed(-16, 8),
    to_signed(-22, 8),
    to_signed(-25, 8),
    to_signed(-25, 8),
    to_signed(-19, 8),
    to_signed(-6, 8),
    to_signed(10, 8),
    to_signed(21, 8),
    to_signed(22, 8),
    to_signed(13, 8),
    to_signed(0, 8),
    to_signed(-13, 8),
    to_signed(-24, 8),
    to_signed(-28, 8),
    to_signed(-24, 8),
    to_signed(-14, 8),
    to_signed(-4, 8),
    to_signed(5, 8),
    to_signed(11, 8),
    to_signed(13, 8),
    to_signed(13, 8),
    to_signed(12, 8),
    to_signed(8, 8),
    to_signed(3, 8),
    to_signed(0, 8),
    to_signed(3, 8),
    to_signed(9, 8),
    to_signed(14, 8),
    to_signed(18, 8),
    to_signed(20, 8),
    to_signed(20, 8),
    to_signed(16, 8),
    to_signed(12, 8),
    to_signed(15, 8),
    to_signed(24, 8),
    to_signed(37, 8),
    to_signed(53, 8),
    to_signed(65, 8),
    to_signed(71, 8),
    to_signed(69, 8),
    to_signed(62, 8),
    to_signed(51, 8),
    to_signed(39, 8),
    to_signed(32, 8),
    to_signed(33, 8),
    to_signed(42, 8),
    to_signed(53, 8),
    to_signed(58, 8),
    to_signed(53, 8),
    to_signed(32, 8),
    to_signed(-4, 8),
    to_signed(-46, 8),
    to_signed(-75, 8),
    to_signed(-80, 8),
    to_signed(-63, 8),
    to_signed(-36, 8),
    to_signed(-10, 8),
    to_signed(7, 8),
    to_signed(8, 8),
    to_signed(-4, 8),
    to_signed(-24, 8),
    to_signed(-44, 8),
    to_signed(-62, 8),
    to_signed(-68, 8),
    to_signed(-58, 8),
    to_signed(-39, 8),
    to_signed(-20, 8),
    to_signed(-6, 8),
    to_signed(6, 8),
    to_signed(14, 8),
    to_signed(16, 8),
    to_signed(17, 8),
    to_signed(19, 8),
    to_signed(23, 8),
    to_signed(23, 8),
    to_signed(15, 8),
    to_signed(1, 8),
    to_signed(-15, 8),
    to_signed(-28, 8),
    to_signed(-37, 8),
    to_signed(-40, 8),
    to_signed(-38, 8),
    to_signed(-31, 8),
    to_signed(-17, 8),
    to_signed(-1, 8),
    to_signed(9, 8),
    to_signed(9, 8),
    to_signed(2, 8),
    to_signed(-7, 8),
    to_signed(-15, 8),
    to_signed(-19, 8),
    to_signed(-19, 8),
    to_signed(-15, 8),
    to_signed(-9, 8),
    to_signed(0, 8),
    to_signed(10, 8),
    to_signed(19, 8),
    to_signed(25, 8),
    to_signed(31, 8),
    to_signed(34, 8),
    to_signed(33, 8),
    to_signed(27, 8),
    to_signed(23, 8),
    to_signed(23, 8),
    to_signed(25, 8),
    to_signed(26, 8),
    to_signed(25, 8),
    to_signed(20, 8),
    to_signed(12, 8),
    to_signed(5, 8),
    to_signed(3, 8),
    to_signed(9, 8),
    to_signed(20, 8),
    to_signed(36, 8),
    to_signed(53, 8),
    to_signed(66, 8),
    to_signed(68, 8),
    to_signed(60, 8),
    to_signed(47, 8),
    to_signed(32, 8),
    to_signed(21, 8),
    to_signed(17, 8),
    to_signed(21, 8),
    to_signed(30, 8),
    to_signed(39, 8),
    to_signed(41, 8),
    to_signed(29, 8),
    to_signed(0, 8),
    to_signed(-41, 8),
    to_signed(-76, 8),
    to_signed(-88, 8),
    to_signed(-74, 8),
    to_signed(-47, 8),
    to_signed(-20, 8),
    to_signed(-2, 8),
    to_signed(1, 8),
    to_signed(-12, 8),
    to_signed(-34, 8),
    to_signed(-57, 8),
    to_signed(-72, 8),
    to_signed(-76, 8),
    to_signed(-64, 8),
    to_signed(-40, 8),
    to_signed(-15, 8),
    to_signed(1, 8),
    to_signed(12, 8),
    to_signed(18, 8),
    to_signed(19, 8),
    to_signed(18, 8),
    to_signed(20, 8),
    to_signed(27, 8),
    to_signed(31, 8),
    to_signed(27, 8),
    to_signed(14, 8),
    to_signed(-1, 8),
    to_signed(-14, 8),
    to_signed(-22, 8),
    to_signed(-24, 8),
    to_signed(-20, 8),
    to_signed(-12, 8),
    to_signed(1, 8),
    to_signed(17, 8),
    to_signed(27, 8),
    to_signed(25, 8),
    to_signed(13, 8),
    to_signed(-2, 8),
    to_signed(-13, 8),
    to_signed(-20, 8),
    to_signed(-22, 8),
    to_signed(-19, 8),
    to_signed(-12, 8),
    to_signed(-3, 8),
    to_signed(8, 8),
    to_signed(17, 8),
    to_signed(23, 8),
    to_signed(26, 8),
    to_signed(28, 8),
    to_signed(26, 8),
    to_signed(20, 8),
    to_signed(13, 8),
    to_signed(10, 8),
    to_signed(12, 8),
    to_signed(14, 8),
    to_signed(14, 8),
    to_signed(12, 8),
    to_signed(7, 8),
    to_signed(3, 8),
    to_signed(2, 8),
    to_signed(7, 8),
    to_signed(16, 8),
    to_signed(26, 8),
    to_signed(37, 8),
    to_signed(47, 8),
    to_signed(48, 8),
    to_signed(39, 8),
    to_signed(27, 8),
    to_signed(18, 8),
    to_signed(15, 8),
    to_signed(18, 8),
    to_signed(27, 8),
    to_signed(39, 8),
    to_signed(50, 8),
    to_signed(53, 8),
    to_signed(43, 8),
    to_signed(17, 8),
    to_signed(-22, 8),
    to_signed(-58, 8),
    to_signed(-74, 8),
    to_signed(-63, 8),
    to_signed(-35, 8),
    to_signed(-7, 8),
    to_signed(12, 8),
    to_signed(16, 8),
    to_signed(3, 8),
    to_signed(-23, 8),
    to_signed(-50, 8),
    to_signed(-66, 8),
    to_signed(-69, 8),
    to_signed(-56, 8),
    to_signed(-33, 8),
    to_signed(-8, 8),
    to_signed(9, 8),
    to_signed(16, 8),
    to_signed(17, 8),
    to_signed(14, 8),
    to_signed(10, 8),
    to_signed(9, 8),
    to_signed(16, 8),
    to_signed(24, 8),
    to_signed(22, 8),
    to_signed(10, 8),
    to_signed(-6, 8),
    to_signed(-21, 8),
    to_signed(-32, 8),
    to_signed(-37, 8),
    to_signed(-36, 8),
    to_signed(-30, 8),
    to_signed(-20, 8),
    to_signed(-6, 8),
    to_signed(5, 8),
    to_signed(4, 8),
    to_signed(-7, 8),
    to_signed(-20, 8),
    to_signed(-30, 8),
    to_signed(-36, 8),
    to_signed(-37, 8),
    to_signed(-31, 8),
    to_signed(-21, 8),
    to_signed(-11, 8),
    to_signed(0, 8),
    to_signed(10, 8),
    to_signed(17, 8),
    to_signed(21, 8),
    to_signed(22, 8),
    to_signed(19, 8),
    to_signed(10, 8),
    to_signed(1, 8),
    to_signed(-3, 8),
    to_signed(0, 8),
    to_signed(6, 8),
    to_signed(10, 8),
    to_signed(10, 8),
    to_signed(8, 8),
    to_signed(6, 8),
    to_signed(5, 8),
    to_signed(7, 8),
    to_signed(14, 8),
    to_signed(23, 8),
    to_signed(33, 8),
    to_signed(42, 8),
    to_signed(46, 8),
    to_signed(40, 8),
    to_signed(28, 8),
    to_signed(17, 8),
    to_signed(14, 8),
    to_signed(18, 8),
    to_signed(30, 8),
    to_signed(46, 8),
    to_signed(60, 8),
    to_signed(64, 8),
    to_signed(54, 8),
    to_signed(28, 8),
    to_signed(-12, 8),
    to_signed(-57, 8),
    to_signed(-87, 8),
    to_signed(-89, 8),
    to_signed(-67, 8),
    to_signed(-36, 8),
    to_signed(-10, 8),
    to_signed(3, 8),
    to_signed(-2, 8),
    to_signed(-22, 8),
    to_signed(-48, 8),
    to_signed(-70, 8),
    to_signed(-79, 8),
    to_signed(-76, 8),
    to_signed(-61, 8),
    to_signed(-40, 8),
    to_signed(-20, 8),
    to_signed(-9, 8),
    to_signed(-2, 8),
    to_signed(3, 8),
    to_signed(6, 8),
    to_signed(7, 8),
    to_signed(14, 8),
    to_signed(23, 8),
    to_signed(25, 8),
    to_signed(16, 8),
    to_signed(-1, 8),
    to_signed(-19, 8),
    to_signed(-34, 8),
    to_signed(-43, 8),
    to_signed(-44, 8),
    to_signed(-40, 8),
    to_signed(-31, 8),
    to_signed(-18, 8),
    to_signed(-3, 8),
    to_signed(3, 8),
    to_signed(-4, 8),
    to_signed(-18, 8),
    to_signed(-29, 8),
    to_signed(-36, 8),
    to_signed(-37, 8),
    to_signed(-33, 8),
    to_signed(-25, 8),
    to_signed(-15, 8),
    to_signed(-6, 8),
    to_signed(3, 8),
    to_signed(11, 8),
    to_signed(17, 8),
    to_signed(20, 8),
    to_signed(22, 8),
    to_signed(19, 8),
    to_signed(13, 8),
    to_signed(9, 8),
    to_signed(10, 8),
    to_signed(14, 8),
    to_signed(15, 8),
    to_signed(10, 8),
    to_signed(2, 8),
    to_signed(-5, 8),
    to_signed(-8, 8),
    to_signed(-6, 8),
    to_signed(0, 8),
    to_signed(9, 8),
    to_signed(20, 8),
    to_signed(31, 8),
    to_signed(37, 8),
    to_signed(33, 8),
    to_signed(22, 8),
    to_signed(10, 8),
    to_signed(4, 8),
    to_signed(6, 8),
    to_signed(15, 8),
    to_signed(30, 8),
    to_signed(47, 8),
    to_signed(58, 8),
    to_signed(57, 8),
    to_signed(42, 8),
    to_signed(12, 8),
    to_signed(-28, 8),
    to_signed(-64, 8),
    to_signed(-78, 8),
    to_signed(-67, 8),
    to_signed(-41, 8),
    to_signed(-14, 8),
    to_signed(5, 8),
    to_signed(8, 8),
    to_signed(-6, 8),
    to_signed(-30, 8),
    to_signed(-51, 8),
    to_signed(-62, 8),
    to_signed(-63, 8),
    to_signed(-52, 8),
    to_signed(-33, 8),
    to_signed(-13, 8),
    to_signed(1, 8),
    to_signed(9, 8),
    to_signed(14, 8),
    to_signed(17, 8),
    to_signed(18, 8),
    to_signed(20, 8),
    to_signed(27, 8),
    to_signed(33, 8),
    to_signed(31, 8),
    to_signed(19, 8),
    to_signed(3, 8),
    to_signed(-13, 8),
    to_signed(-26, 8),
    to_signed(-34, 8),
    to_signed(-37, 8),
    to_signed(-34, 8),
    to_signed(-25, 8),
    to_signed(-11, 8),
    to_signed(-2, 8),
    to_signed(-6, 8),
    to_signed(-21, 8),
    to_signed(-36, 8),
    to_signed(-46, 8),
    to_signed(-49, 8),
    to_signed(-44, 8),
    to_signed(-34, 8),
    to_signed(-23, 8),
    to_signed(-12, 8),
    to_signed(-1, 8),
    to_signed(7, 8),
    to_signed(15, 8),
    to_signed(21, 8),
    to_signed(25, 8),
    to_signed(25, 8),
    to_signed(20, 8),
    to_signed(14, 8),
    to_signed(14, 8),
    to_signed(20, 8),
    to_signed(27, 8),
    to_signed(31, 8),
    to_signed(31, 8),
    to_signed(29, 8),
    to_signed(25, 8),
    to_signed(21, 8),
    to_signed(18, 8),
    to_signed(19, 8),
    to_signed(25, 8),
    to_signed(35, 8),
    to_signed(47, 8),
    to_signed(52, 8),
    to_signed(49, 8),
    to_signed(43, 8),
    to_signed(39, 8),
    to_signed(39, 8),
    to_signed(44, 8),
    to_signed(53, 8),
    to_signed(64, 8),
    to_signed(75, 8),
    to_signed(77, 8),
    to_signed(67, 8),
    to_signed(43, 8),
    to_signed(5, 8),
    to_signed(-35, 8),
    to_signed(-63, 8),
    to_signed(-68, 8),
    to_signed(-50, 8),
    to_signed(-26, 8),
    to_signed(-6, 8),
    to_signed(3, 8),
    to_signed(-2, 8),
    to_signed(-21, 8),
    to_signed(-45, 8),
    to_signed(-63, 8),
    to_signed(-72, 8),
    to_signed(-71, 8),
    to_signed(-60, 8),
    to_signed(-43, 8),
    to_signed(-27, 8),
    to_signed(-17, 8),
    to_signed(-10, 8),
    to_signed(-3, 8),
    to_signed(2, 8),
    to_signed(7, 8),
    to_signed(13, 8),
    to_signed(21, 8),
    to_signed(23, 8),
    to_signed(16, 8),
    to_signed(2, 8),
    to_signed(-15, 8),
    to_signed(-31, 8),
    to_signed(-43, 8),
    to_signed(-50, 8),
    to_signed(-50, 8),
    to_signed(-39, 8),
    to_signed(-19, 8),
    to_signed(0, 8),
    to_signed(8, 8),
    to_signed(3, 8),
    to_signed(-10, 8),
    to_signed(-24, 8),
    to_signed(-34, 8),
    to_signed(-36, 8),
    to_signed(-30, 8),
    to_signed(-19, 8),
    to_signed(-5, 8),
    to_signed(8, 8),
    to_signed(21, 8),
    to_signed(30, 8),
    to_signed(37, 8),
    to_signed(43, 8),
    to_signed(46, 8),
    to_signed(42, 8),
    to_signed(35, 8),
    to_signed(30, 8),
    to_signed(29, 8),
    to_signed(33, 8),
    to_signed(36, 8),
    to_signed(37, 8),
    to_signed(35, 8),
    to_signed(30, 8),
    to_signed(24, 8),
    to_signed(18, 8),
    to_signed(16, 8),
    to_signed(19, 8),
    to_signed(26, 8),
    to_signed(35, 8),
    to_signed(41, 8),
    to_signed(40, 8),
    to_signed(32, 8),
    to_signed(25, 8),
    to_signed(23, 8),
    to_signed(25, 8),
    to_signed(31, 8),
    to_signed(40, 8),
    to_signed(49, 8),
    to_signed(55, 8),
    to_signed(52, 8),
    to_signed(35, 8),
    to_signed(4, 8),
    to_signed(-37, 8),
    to_signed(-71, 8),
    to_signed(-84, 8),
    to_signed(-74, 8),
    to_signed(-51, 8),
    to_signed(-29, 8),
    to_signed(-16, 8),
    to_signed(-14, 8),
    to_signed(-25, 8),
    to_signed(-44, 8),
    to_signed(-64, 8),
    to_signed(-75, 8),
    to_signed(-75, 8),
    to_signed(-65, 8),
    to_signed(-49, 8),
    to_signed(-30, 8),
    to_signed(-14, 8),
    to_signed(-3, 8),
    to_signed(5, 8),
    to_signed(10, 8),
    to_signed(14, 8),
    to_signed(20, 8),
    to_signed(29, 8),
    to_signed(36, 8),
    to_signed(34, 8),
    to_signed(25, 8),
    to_signed(10, 8),
    to_signed(-7, 8),
    to_signed(-24, 8),
    to_signed(-37, 8),
    to_signed(-42, 8),
    to_signed(-36, 8),
    to_signed(-18, 8),
    to_signed(5, 8),
    to_signed(20, 8),
    to_signed(19, 8),
    to_signed(8, 8),
    to_signed(-7, 8),
    to_signed(-21, 8),
    to_signed(-30, 8),
    to_signed(-29, 8),
    to_signed(-19, 8),
    to_signed(-6, 8),
    to_signed(6, 8),
    to_signed(15, 8),
    to_signed(20, 8),
    to_signed(24, 8),
    to_signed(28, 8),
    to_signed(33, 8),
    to_signed(33, 8),
    to_signed(27, 8),
    to_signed(20, 8),
    to_signed(15, 8),
    to_signed(14, 8),
    to_signed(14, 8),
    to_signed(15, 8),
    to_signed(14, 8),
    to_signed(11, 8),
    to_signed(6, 8),
    to_signed(1, 8),
    to_signed(0, 8),
    to_signed(3, 8),
    to_signed(12, 8),
    to_signed(22, 8),
    to_signed(32, 8),
    to_signed(35, 8),
    to_signed(33, 8),
    to_signed(27, 8),
    to_signed(23, 8),
    to_signed(23, 8),
    to_signed(26, 8),
    to_signed(32, 8),
    to_signed(40, 8),
    to_signed(49, 8),
    to_signed(53, 8),
    to_signed(46, 8),
    to_signed(24, 8),
    to_signed(-12, 8),
    to_signed(-51, 8),
    to_signed(-77, 8),
    to_signed(-78, 8),
    to_signed(-60, 8),
    to_signed(-37, 8),
    to_signed(-18, 8),
    to_signed(-8, 8),
    to_signed(-10, 8),
    to_signed(-24, 8),
    to_signed(-43, 8),
    to_signed(-57, 8),
    to_signed(-62, 8),
    to_signed(-56, 8),
    to_signed(-41, 8),
    to_signed(-23, 8),
    to_signed(-6, 8),
    to_signed(6, 8),
    to_signed(14, 8),
    to_signed(20, 8),
    to_signed(22, 8),
    to_signed(23, 8),
    to_signed(28, 8),
    to_signed(33, 8),
    to_signed(33, 8),
    to_signed(24, 8),
    to_signed(10, 8),
    to_signed(-5, 8),
    to_signed(-20, 8),
    to_signed(-33, 8),
    to_signed(-43, 8),
    to_signed(-45, 8),
    to_signed(-37, 8),
    to_signed(-22, 8),
    to_signed(-8, 8),
    to_signed(-3, 8),
    to_signed(-8, 8),
    to_signed(-18, 8),
    to_signed(-27, 8),
    to_signed(-35, 8),
    to_signed(-40, 8),
    to_signed(-37, 8),
    to_signed(-27, 8),
    to_signed(-15, 8),
    to_signed(-4, 8),
    to_signed(4, 8),
    to_signed(10, 8),
    to_signed(15, 8),
    to_signed(21, 8),
    to_signed(24, 8),
    to_signed(21, 8),
    to_signed(13, 8),
    to_signed(8, 8),
    to_signed(9, 8),
    to_signed(10, 8),
    to_signed(12, 8),
    to_signed(12, 8),
    to_signed(10, 8),
    to_signed(7, 8),
    to_signed(2, 8),
    to_signed(-2, 8),
    to_signed(-4, 8),
    to_signed(-1, 8),
    to_signed(6, 8),
    to_signed(15, 8),
    to_signed(23, 8),
    to_signed(27, 8),
    to_signed(29, 8),
    to_signed(30, 8),
    to_signed(30, 8),
    to_signed(30, 8),
    to_signed(30, 8),
    to_signed(31, 8),
    to_signed(36, 8),
    to_signed(45, 8),
    to_signed(50, 8),
    to_signed(44, 8),
    to_signed(24, 8),
    to_signed(-8, 8),
    to_signed(-41, 8),
    to_signed(-60, 8),
    to_signed(-59, 8),
    to_signed(-47, 8),
    to_signed(-33, 8),
    to_signed(-23, 8),
    to_signed(-19, 8),
    to_signed(-25, 8),
    to_signed(-38, 8),
    to_signed(-50, 8),
    to_signed(-55, 8),
    to_signed(-55, 8),
    to_signed(-49, 8),
    to_signed(-37, 8),
    to_signed(-25, 8),
    to_signed(-17, 8),
    to_signed(-10, 8),
    to_signed(-3, 8),
    to_signed(4, 8),
    to_signed(11, 8),
    to_signed(20, 8),
    to_signed(31, 8),
    to_signed(38, 8),
    to_signed(36, 8),
    to_signed(24, 8),
    to_signed(7, 8),
    to_signed(-10, 8),
    to_signed(-26, 8),
    to_signed(-38, 8),
    to_signed(-44, 8),
    to_signed(-40, 8),
    to_signed(-27, 8),
    to_signed(-12, 8),
    to_signed(-2, 8),
    to_signed(-1, 8),
    to_signed(-8, 8),
    to_signed(-19, 8),
    to_signed(-28, 8),
    to_signed(-34, 8),
    to_signed(-34, 8),
    to_signed(-28, 8),
    to_signed(-16, 8),
    to_signed(-5, 8),
    to_signed(2, 8),
    to_signed(6, 8),
    to_signed(10, 8),
    to_signed(14, 8),
    to_signed(18, 8),
    to_signed(18, 8),
    to_signed(13, 8),
    to_signed(7, 8),
    to_signed(7, 8),
    to_signed(13, 8),
    to_signed(19, 8),
    to_signed(22, 8),
    to_signed(20, 8),
    to_signed(15, 8),
    to_signed(7, 8),
    to_signed(0, 8),
    to_signed(-5, 8),
    to_signed(-4, 8),
    to_signed(2, 8),
    to_signed(15, 8),
    to_signed(29, 8),
    to_signed(38, 8),
    to_signed(42, 8),
    to_signed(44, 8),
    to_signed(44, 8),
    to_signed(43, 8),
    to_signed(41, 8),
    to_signed(41, 8),
    to_signed(45, 8),
    to_signed(54, 8),
    to_signed(64, 8),
    to_signed(67, 8),
    to_signed(55, 8),
    to_signed(28, 8),
    to_signed(-7, 8),
    to_signed(-38, 8),
    to_signed(-51, 8),
    to_signed(-45, 8),
    to_signed(-29, 8),
    to_signed(-13, 8),
    to_signed(0, 8),
    to_signed(3, 8),
    to_signed(-6, 8),
    to_signed(-23, 8),
    to_signed(-37, 8),
    to_signed(-45, 8),
    to_signed(-50, 8),
    to_signed(-47, 8),
    to_signed(-36, 8),
    to_signed(-26, 8),
    to_signed(-20, 8),
    to_signed(-15, 8),
    to_signed(-6, 8),
    to_signed(2, 8),
    to_signed(11, 8),
    to_signed(25, 8),
    to_signed(38, 8),
    to_signed(43, 8),
    to_signed(33, 8),
    to_signed(14, 8),
    to_signed(-9, 8),
    to_signed(-30, 8),
    to_signed(-45, 8),
    to_signed(-54, 8),
    to_signed(-54, 8),
    to_signed(-44, 8),
    to_signed(-29, 8),
    to_signed(-13, 8),
    to_signed(-3, 8),
    to_signed(1, 8),
    to_signed(-3, 8),
    to_signed(-12, 8),
    to_signed(-19, 8),
    to_signed(-23, 8),
    to_signed(-26, 8),
    to_signed(-25, 8),
    to_signed(-19, 8),
    to_signed(-10, 8),
    to_signed(-2, 8),
    to_signed(8, 8),
    to_signed(21, 8),
    to_signed(34, 8),
    to_signed(43, 8),
    to_signed(44, 8),
    to_signed(39, 8),
    to_signed(34, 8),
    to_signed(33, 8),
    to_signed(35, 8),
    to_signed(36, 8),
    to_signed(32, 8),
    to_signed(26, 8),
    to_signed(19, 8),
    to_signed(14, 8),
    to_signed(11, 8),
    to_signed(12, 8),
    to_signed(17, 8),
    to_signed(26, 8),
    to_signed(38, 8),
    to_signed(46, 8),
    to_signed(47, 8),
    to_signed(42, 8),
    to_signed(37, 8),
    to_signed(32, 8),
    to_signed(27, 8),
    to_signed(25, 8),
    to_signed(26, 8),
    to_signed(29, 8),
    to_signed(36, 8),
    to_signed(41, 8),
    to_signed(36, 8),
    to_signed(15, 8),
    to_signed(-17, 8),
    to_signed(-48, 8),
    to_signed(-67, 8),
    to_signed(-67, 8),
    to_signed(-54, 8),
    to_signed(-39, 8),
    to_signed(-28, 8),
    to_signed(-26, 8),
    to_signed(-33, 8),
    to_signed(-49, 8),
    to_signed(-66, 8),
    to_signed(-73, 8),
    to_signed(-73, 8),
    to_signed(-65, 8),
    to_signed(-52, 8),
    to_signed(-36, 8),
    to_signed(-25, 8),
    to_signed(-21, 8),
    to_signed(-18, 8),
    to_signed(-13, 8),
    to_signed(-8, 8),
    to_signed(3, 8),
    to_signed(20, 8),
    to_signed(36, 8),
    to_signed(41, 8),
    to_signed(32, 8),
    to_signed(15, 8),
    to_signed(-3, 8),
    to_signed(-19, 8),
    to_signed(-31, 8),
    to_signed(-36, 8),
    to_signed(-31, 8),
    to_signed(-17, 8),
    to_signed(-1, 8),
    to_signed(10, 8),
    to_signed(13, 8),
    to_signed(6, 8),
    to_signed(-6, 8),
    to_signed(-18, 8),
    to_signed(-24, 8),
    to_signed(-22, 8),
    to_signed(-17, 8),
    to_signed(-9, 8),
    to_signed(-2, 8),
    to_signed(5, 8),
    to_signed(10, 8),
    to_signed(17, 8),
    to_signed(25, 8),
    to_signed(30, 8),
    to_signed(30, 8),
    to_signed(24, 8),
    to_signed(16, 8),
    to_signed(13, 8),
    to_signed(15, 8),
    to_signed(19, 8),
    to_signed(21, 8),
    to_signed(18, 8),
    to_signed(12, 8),
    to_signed(2, 8),
    to_signed(-7, 8),
    to_signed(-12, 8),
    to_signed(-12, 8),
    to_signed(-6, 8),
    to_signed(5, 8),
    to_signed(18, 8),
    to_signed(25, 8),
    to_signed(24, 8),
    to_signed(17, 8),
    to_signed(10, 8),
    to_signed(7, 8),
    to_signed(9, 8),
    to_signed(13, 8),
    to_signed(19, 8),
    to_signed(27, 8),
    to_signed(35, 8),
    to_signed(37, 8),
    to_signed(24, 8),
    to_signed(-3, 8),
    to_signed(-37, 8),
    to_signed(-66, 8),
    to_signed(-77, 8),
    to_signed(-69, 8),
    to_signed(-50, 8),
    to_signed(-31, 8),
    to_signed(-16, 8),
    to_signed(-11, 8),
    to_signed(-19, 8),
    to_signed(-36, 8),
    to_signed(-53, 8),
    to_signed(-61, 8),
    to_signed(-58, 8),
    to_signed(-48, 8),
    to_signed(-33, 8),
    to_signed(-19, 8),
    to_signed(-11, 8),
    to_signed(-7, 8),
    to_signed(-4, 8),
    to_signed(0, 8),
    to_signed(9, 8),
    to_signed(24, 8),
    to_signed(40, 8),
    to_signed(51, 8),
    to_signed(47, 8),
    to_signed(30, 8),
    to_signed(9, 8),
    to_signed(-8, 8),
    to_signed(-20, 8),
    to_signed(-28, 8),
    to_signed(-27, 8),
    to_signed(-16, 8),
    to_signed(0, 8),
    to_signed(14, 8),
    to_signed(21, 8),
    to_signed(19, 8),
    to_signed(9, 8),
    to_signed(-3, 8),
    to_signed(-14, 8),
    to_signed(-19, 8),
    to_signed(-19, 8),
    to_signed(-14, 8),
    to_signed(-8, 8),
    to_signed(-2, 8),
    to_signed(4, 8),
    to_signed(10, 8),
    to_signed(17, 8),
    to_signed(22, 8),
    to_signed(25, 8),
    to_signed(23, 8),
    to_signed(18, 8),
    to_signed(15, 8),
    to_signed(15, 8),
    to_signed(17, 8),
    to_signed(18, 8),
    to_signed(17, 8),
    to_signed(14, 8),
    to_signed(7, 8),
    to_signed(0, 8),
    to_signed(-6, 8),
    to_signed(-8, 8),
    to_signed(-6, 8),
    to_signed(3, 8),
    to_signed(17, 8),
    to_signed(29, 8),
    to_signed(36, 8),
    to_signed(35, 8),
    to_signed(27, 8),
    to_signed(17, 8),
    to_signed(14, 8),
    to_signed(17, 8),
    to_signed(23, 8),
    to_signed(29, 8),
    to_signed(37, 8),
    to_signed(42, 8),
    to_signed(38, 8),
    to_signed(20, 8),
    to_signed(-9, 8),
    to_signed(-38, 8),
    to_signed(-56, 8),
    to_signed(-57, 8),
    to_signed(-45, 8),
    to_signed(-28, 8),
    to_signed(-15, 8),
    to_signed(-9, 8),
    to_signed(-12, 8),
    to_signed(-22, 8),
    to_signed(-36, 8),
    to_signed(-47, 8),
    to_signed(-49, 8),
    to_signed(-40, 8),
    to_signed(-25, 8),
    to_signed(-12, 8),
    to_signed(-1, 8),
    to_signed(9, 8),
    to_signed(16, 8),
    to_signed(19, 8),
    to_signed(23, 8),
    to_signed(33, 8),
    to_signed(46, 8),
    to_signed(57, 8),
    to_signed(60, 8),
    to_signed(51, 8),
    to_signed(31, 8),
    to_signed(8, 8),
    to_signed(-9, 8),
    to_signed(-22, 8),
    to_signed(-30, 8),
    to_signed(-28, 8),
    to_signed(-17, 8),
    to_signed(-2, 8),
    to_signed(8, 8),
    to_signed(10, 8),
    to_signed(1, 8),
    to_signed(-13, 8),
    to_signed(-27, 8),
    to_signed(-36, 8),
    to_signed(-40, 8),
    to_signed(-37, 8),
    to_signed(-25, 8),
    to_signed(-13, 8),
    to_signed(-3, 8),
    to_signed(8, 8),
    to_signed(17, 8),
    to_signed(23, 8),
    to_signed(25, 8),
    to_signed(24, 8),
    to_signed(19, 8),
    to_signed(11, 8),
    to_signed(6, 8),
    to_signed(7, 8),
    to_signed(7, 8),
    to_signed(5, 8),
    to_signed(2, 8),
    to_signed(-4, 8),
    to_signed(-12, 8),
    to_signed(-18, 8),
    to_signed(-20, 8),
    to_signed(-20, 8),
    to_signed(-14, 8),
    to_signed(-1, 8),
    to_signed(13, 8),
    to_signed(22, 8),
    to_signed(26, 8),
    to_signed(25, 8),
    to_signed(17, 8),
    to_signed(10, 8),
    to_signed(13, 8),
    to_signed(24, 8),
    to_signed(35, 8),
    to_signed(45, 8),
    to_signed(54, 8),
    to_signed(57, 8),
    to_signed(47, 8),
    to_signed(23, 8),
    to_signed(-10, 8),
    to_signed(-40, 8),
    to_signed(-54, 8),
    to_signed(-49, 8),
    to_signed(-32, 8),
    to_signed(-15, 8),
    to_signed(-4, 8),
    to_signed(-3, 8),
    to_signed(-14, 8),
    to_signed(-29, 8),
    to_signed(-44, 8),
    to_signed(-55, 8),
    to_signed(-57, 8),
    to_signed(-47, 8),
    to_signed(-34, 8),
    to_signed(-25, 8),
    to_signed(-18, 8),
    to_signed(-11, 8),
    to_signed(-4, 8),
    to_signed(0, 8),
    to_signed(6, 8),
    to_signed(18, 8),
    to_signed(31, 8),
    to_signed(38, 8),
    to_signed(36, 8),
    to_signed(23, 8),
    to_signed(4, 8),
    to_signed(-12, 8),
    to_signed(-22, 8),
    to_signed(-29, 8),
    to_signed(-30, 8),
    to_signed(-23, 8),
    to_signed(-11, 8),
    to_signed(4, 8),
    to_signed(15, 8),
    to_signed(18, 8),
    to_signed(10, 8),
    to_signed(-4, 8),
    to_signed(-15, 8),
    to_signed(-25, 8),
    to_signed(-33, 8),
    to_signed(-30, 8),
    to_signed(-17, 8),
    to_signed(-2, 8),
    to_signed(11, 8),
    to_signed(25, 8),
    to_signed(38, 8),
    to_signed(47, 8),
    to_signed(52, 8),
    to_signed(50, 8),
    to_signed(42, 8),
    to_signed(33, 8),
    to_signed(28, 8),
    to_signed(28, 8),
    to_signed(28, 8),
    to_signed(28, 8),
    to_signed(27, 8),
    to_signed(24, 8),
    to_signed(19, 8),
    to_signed(16, 8),
    to_signed(15, 8),
    to_signed(14, 8),
    to_signed(19, 8),
    to_signed(28, 8),
    to_signed(34, 8),
    to_signed(34, 8),
    to_signed(29, 8),
    to_signed(20, 8),
    to_signed(8, 8),
    to_signed(1, 8),
    to_signed(8, 8),
    to_signed(25, 8),
    to_signed(44, 8),
    to_signed(59, 8),
    to_signed(67, 8),
    to_signed(63, 8),
    to_signed(44, 8),
    to_signed(11, 8),
    to_signed(-28, 8),
    to_signed(-61, 8),
    to_signed(-75, 8),
    to_signed(-67, 8),
    to_signed(-48, 8),
    to_signed(-29, 8),
    to_signed(-16, 8),
    to_signed(-11, 8),
    to_signed(-15, 8),
    to_signed(-24, 8),
    to_signed(-36, 8),
    to_signed(-46, 8),
    to_signed(-49, 8),
    to_signed(-44, 8),
    to_signed(-35, 8),
    to_signed(-29, 8),
    to_signed(-23, 8),
    to_signed(-13, 8),
    to_signed(-2, 8),
    to_signed(12, 8),
    to_signed(28, 8),
    to_signed(48, 8),
    to_signed(63, 8),
    to_signed(68, 8),
    to_signed(57, 8),
    to_signed(32, 8),
    to_signed(4, 8),
    to_signed(-16, 8),
    to_signed(-27, 8),
    to_signed(-33, 8),
    to_signed(-30, 8),
    to_signed(-19, 8),
    to_signed(-4, 8),
    to_signed(8, 8),
    to_signed(15, 8),
    to_signed(13, 8),
    to_signed(4, 8),
    to_signed(-7, 8),
    to_signed(-16, 8),
    to_signed(-25, 8),
    to_signed(-33, 8),
    to_signed(-34, 8),
    to_signed(-25, 8),
    to_signed(-13, 8),
    to_signed(-2, 8),
    to_signed(10, 8),
    to_signed(22, 8),
    to_signed(32, 8),
    to_signed(35, 8),
    to_signed(29, 8),
    to_signed(17, 8),
    to_signed(8, 8),
    to_signed(6, 8),
    to_signed(6, 8),
    to_signed(5, 8),
    to_signed(4, 8),
    to_signed(2, 8),
    to_signed(-4, 8),
    to_signed(-12, 8),
    to_signed(-15, 8),
    to_signed(-15, 8),
    to_signed(-11, 8),
    to_signed(-2, 8),
    to_signed(13, 8),
    to_signed(26, 8),
    to_signed(31, 8),
    to_signed(30, 8),
    to_signed(22, 8),
    to_signed(10, 8),
    to_signed(2, 8),
    to_signed(6, 8),
    to_signed(19, 8),
    to_signed(36, 8),
    to_signed(51, 8),
    to_signed(60, 8),
    to_signed(58, 8),
    to_signed(43, 8),
    to_signed(14, 8),
    to_signed(-23, 8),
    to_signed(-54, 8),
    to_signed(-64, 8),
    to_signed(-54, 8),
    to_signed(-37, 8),
    to_signed(-22, 8),
    to_signed(-11, 8),
    to_signed(-8, 8),
    to_signed(-13, 8),
    to_signed(-23, 8),
    to_signed(-32, 8),
    to_signed(-38, 8),
    to_signed(-38, 8),
    to_signed(-33, 8),
    to_signed(-26, 8),
    to_signed(-22, 8),
    to_signed(-20, 8),
    to_signed(-16, 8),
    to_signed(-8, 8),
    to_signed(5, 8),
    to_signed(21, 8),
    to_signed(38, 8),
    to_signed(50, 8),
    to_signed(51, 8),
    to_signed(35, 8),
    to_signed(9, 8),
    to_signed(-17, 8),
    to_signed(-35, 8),
    to_signed(-46, 8),
    to_signed(-50, 8),
    to_signed(-46, 8),
    to_signed(-33, 8),
    to_signed(-19, 8),
    to_signed(-9, 8),
    to_signed(-5, 8),
    to_signed(-11, 8),
    to_signed(-24, 8),
    to_signed(-37, 8),
    to_signed(-47, 8),
    to_signed(-54, 8),
    to_signed(-56, 8),
    to_signed(-51, 8),
    to_signed(-39, 8),
    to_signed(-26, 8),
    to_signed(-14, 8),
    to_signed(-2, 8),
    to_signed(8, 8),
    to_signed(16, 8),
    to_signed(17, 8),
    to_signed(11, 8),
    to_signed(-1, 8),
    to_signed(-7, 8),
    to_signed(-6, 8),
    to_signed(-1, 8),
    to_signed(2, 8),
    to_signed(5, 8),
    to_signed(7, 8),
    to_signed(6, 8),
    to_signed(-1, 8),
    to_signed(-9, 8),
    to_signed(-13, 8),
    to_signed(-10, 8),
    to_signed(1, 8),
    to_signed(16, 8),
    to_signed(31, 8),
    to_signed(38, 8),
    to_signed(36, 8),
    to_signed(29, 8),
    to_signed(19, 8),
    to_signed(12, 8),
    to_signed(13, 8),
    to_signed(22, 8),
    to_signed(34, 8),
    to_signed(47, 8),
    to_signed(53, 8),
    to_signed(49, 8),
    to_signed(32, 8),
    to_signed(2, 8),
    to_signed(-38, 8),
    to_signed(-74, 8),
    to_signed(-89, 8),
    to_signed(-81, 8),
    to_signed(-63, 8),
    to_signed(-45, 8),
    to_signed(-31, 8),
    to_signed(-23, 8),
    to_signed(-27, 8),
    to_signed(-39, 8),
    to_signed(-51, 8),
    to_signed(-59, 8),
    to_signed(-63, 8),
    to_signed(-60, 8),
    to_signed(-50, 8),
    to_signed(-39, 8),
    to_signed(-31, 8),
    to_signed(-24, 8),
    to_signed(-12, 8),
    to_signed(2, 8),
    to_signed(19, 8),
    to_signed(36, 8),
    to_signed(48, 8),
    to_signed(47, 8),
    to_signed(32, 8),
    to_signed(8, 8),
    to_signed(-15, 8),
    to_signed(-29, 8),
    to_signed(-38, 8),
    to_signed(-40, 8),
    to_signed(-35, 8),
    to_signed(-23, 8),
    to_signed(-9, 8),
    to_signed(2, 8),
    to_signed(8, 8),
    to_signed(7, 8),
    to_signed(-2, 8),
    to_signed(-12, 8),
    to_signed(-21, 8),
    to_signed(-28, 8),
    to_signed(-33, 8),
    to_signed(-31, 8),
    to_signed(-21, 8),
    to_signed(-7, 8),
    to_signed(6, 8),
    to_signed(16, 8),
    to_signed(26, 8),
    to_signed(32, 8),
    to_signed(32, 8),
    to_signed(23, 8),
    to_signed(11, 8),
    to_signed(2, 8),
    to_signed(1, 8),
    to_signed(4, 8),
    to_signed(6, 8),
    to_signed(6, 8),
    to_signed(7, 8),
    to_signed(6, 8),
    to_signed(2, 8),
    to_signed(-7, 8),
    to_signed(-16, 8),
    to_signed(-17, 8),
    to_signed(-9, 8),
    to_signed(6, 8),
    to_signed(20, 8),
    to_signed(29, 8),
    to_signed(31, 8),
    to_signed(28, 8),
    to_signed(23, 8),
    to_signed(21, 8),
    to_signed(25, 8),
    to_signed(32, 8),
    to_signed(43, 8),
    to_signed(55, 8),
    to_signed(63, 8),
    to_signed(62, 8),
    to_signed(49, 8),
    to_signed(23, 8),
    to_signed(-16, 8),
    to_signed(-53, 8),
    to_signed(-71, 8),
    to_signed(-64, 8),
    to_signed(-45, 8),
    to_signed(-26, 8),
    to_signed(-10, 8),
    to_signed(3, 8),
    to_signed(5, 8),
    to_signed(-6, 8),
    to_signed(-25, 8),
    to_signed(-42, 8),
    to_signed(-55, 8),
    to_signed(-57, 8),
    to_signed(-50, 8),
    to_signed(-36, 8),
    to_signed(-22, 8),
    to_signed(-8, 8),
    to_signed(7, 8),
    to_signed(24, 8),
    to_signed(39, 8),
    to_signed(52, 8),
    to_signed(60, 8),
    to_signed(58, 8),
    to_signed(42, 8),
    to_signed(17, 8),
    to_signed(-9, 8),
    to_signed(-29, 8),
    to_signed(-39, 8),
    to_signed(-42, 8),
    to_signed(-36, 8),
    to_signed(-23, 8),
    to_signed(-8, 8),
    to_signed(4, 8),
    to_signed(10, 8),
    to_signed(8, 8),
    to_signed(-2, 8),
    to_signed(-15, 8),
    to_signed(-28, 8),
    to_signed(-36, 8),
    to_signed(-39, 8),
    to_signed(-36, 8),
    to_signed(-26, 8),
    to_signed(-10, 8),
    to_signed(8, 8),
    to_signed(25, 8),
    to_signed(38, 8),
    to_signed(46, 8),
    to_signed(46, 8),
    to_signed(38, 8),
    to_signed(27, 8),
    to_signed(19, 8),
    to_signed(19, 8),
    to_signed(23, 8),
    to_signed(25, 8),
    to_signed(26, 8),
    to_signed(27, 8),
    to_signed(26, 8),
    to_signed(22, 8),
    to_signed(14, 8),
    to_signed(7, 8),
    to_signed(5, 8),
    to_signed(12, 8),
    to_signed(27, 8),
    to_signed(42, 8),
    to_signed(52, 8),
    to_signed(57, 8),
    to_signed(57, 8),
    to_signed(50, 8),
    to_signed(40, 8),
    to_signed(34, 8),
    to_signed(34, 8),
    to_signed(39, 8),
    to_signed(51, 8),
    to_signed(64, 8),
    to_signed(72, 8),
    to_signed(66, 8),
    to_signed(44, 8),
    to_signed(6, 8),
    to_signed(-36, 8),
    to_signed(-63, 8),
    to_signed(-67, 8),
    to_signed(-54, 8),
    to_signed(-38, 8),
    to_signed(-23, 8),
    to_signed(-12, 8),
    to_signed(-7, 8),
    to_signed(-13, 8),
    to_signed(-26, 8),
    to_signed(-41, 8),
    to_signed(-54, 8),
    to_signed(-60, 8),
    to_signed(-58, 8),
    to_signed(-50, 8),
    to_signed(-38, 8),
    to_signed(-25, 8),
    to_signed(-8, 8),
    to_signed(10, 8),
    to_signed(29, 8),
    to_signed(45, 8),
    to_signed(53, 8),
    to_signed(49, 8),
    to_signed(34, 8),
    to_signed(13, 8),
    to_signed(-8, 8),
    to_signed(-23, 8),
    to_signed(-30, 8),
    to_signed(-30, 8),
    to_signed(-25, 8),
    to_signed(-13, 8),
    to_signed(2, 8),
    to_signed(12, 8),
    to_signed(15, 8),
    to_signed(11, 8),
    to_signed(0, 8),
    to_signed(-13, 8),
    to_signed(-24, 8),
    to_signed(-32, 8),
    to_signed(-33, 8),
    to_signed(-26, 8),
    to_signed(-14, 8),
    to_signed(1, 8),
    to_signed(18, 8),
    to_signed(34, 8),
    to_signed(45, 8),
    to_signed(50, 8),
    to_signed(46, 8),
    to_signed(35, 8),
    to_signed(21, 8),
    to_signed(12, 8),
    to_signed(12, 8),
    to_signed(17, 8),
    to_signed(24, 8),
    to_signed(28, 8),
    to_signed(30, 8),
    to_signed(28, 8),
    to_signed(21, 8),
    to_signed(8, 8),
    to_signed(-6, 8),
    to_signed(-14, 8),
    to_signed(-9, 8),
    to_signed(6, 8),
    to_signed(23, 8),
    to_signed(36, 8),
    to_signed(43, 8),
    to_signed(42, 8),
    to_signed(36, 8),
    to_signed(29, 8),
    to_signed(23, 8),
    to_signed(20, 8),
    to_signed(22, 8),
    to_signed(31, 8),
    to_signed(45, 8),
    to_signed(53, 8),
    to_signed(51, 8),
    to_signed(32, 8),
    to_signed(-2, 8),
    to_signed(-41, 8),
    to_signed(-70, 8),
    to_signed(-79, 8),
    to_signed(-70, 8),
    to_signed(-53, 8),
    to_signed(-35, 8),
    to_signed(-21, 8),
    to_signed(-15, 8),
    to_signed(-20, 8),
    to_signed(-33, 8),
    to_signed(-49, 8),
    to_signed(-62, 8),
    to_signed(-67, 8),
    to_signed(-65, 8),
    to_signed(-58, 8),
    to_signed(-46, 8),
    to_signed(-29, 8),
    to_signed(-9, 8),
    to_signed(10, 8),
    to_signed(26, 8),
    to_signed(38, 8),
    to_signed(45, 8),
    to_signed(41, 8),
    to_signed(25, 8),
    to_signed(3, 8),
    to_signed(-17, 8),
    to_signed(-30, 8),
    to_signed(-34, 8),
    to_signed(-31, 8),
    to_signed(-24, 8),
    to_signed(-13, 8),
    to_signed(0, 8),
    to_signed(11, 8),
    to_signed(16, 8),
    to_signed(13, 8),
    to_signed(3, 8),
    to_signed(-11, 8),
    to_signed(-24, 8),
    to_signed(-33, 8),
    to_signed(-36, 8),
    to_signed(-32, 8),
    to_signed(-20, 8),
    to_signed(-4, 8),
    to_signed(14, 8),
    to_signed(30, 8),
    to_signed(40, 8),
    to_signed(42, 8),
    to_signed(34, 8),
    to_signed(20, 8),
    to_signed(6, 8),
    to_signed(-3, 8),
    to_signed(-6, 8),
    to_signed(-3, 8),
    to_signed(4, 8),
    to_signed(14, 8),
    to_signed(21, 8),
    to_signed(21, 8),
    to_signed(14, 8),
    to_signed(2, 8),
    to_signed(-13, 8),
    to_signed(-23, 8),
    to_signed(-21, 8),
    to_signed(-9, 8),
    to_signed(6, 8),
    to_signed(18, 8),
    to_signed(25, 8),
    to_signed(24, 8),
    to_signed(17, 8),
    to_signed(12, 8),
    to_signed(11, 8),
    to_signed(13, 8),
    to_signed(19, 8),
    to_signed(30, 8),
    to_signed(43, 8),
    to_signed(51, 8),
    to_signed(48, 8),
    to_signed(30, 8),
    to_signed(-4, 8),
    to_signed(-45, 8),
    to_signed(-75, 8),
    to_signed(-83, 8),
    to_signed(-71, 8),
    to_signed(-49, 8),
    to_signed(-25, 8),
    to_signed(-5, 8),
    to_signed(5, 8),
    to_signed(2, 8),
    to_signed(-15, 8),
    to_signed(-38, 8),
    to_signed(-59, 8),
    to_signed(-71, 8),
    to_signed(-69, 8),
    to_signed(-57, 8),
    to_signed(-39, 8),
    to_signed(-18, 8),
    to_signed(6, 8),
    to_signed(28, 8),
    to_signed(44, 8),
    to_signed(53, 8),
    to_signed(58, 8),
    to_signed(58, 8),
    to_signed(49, 8),
    to_signed(30, 8),
    to_signed(9, 8),
    to_signed(-7, 8),
    to_signed(-18, 8),
    to_signed(-24, 8),
    to_signed(-22, 8),
    to_signed(-13, 8),
    to_signed(0, 8),
    to_signed(11, 8),
    to_signed(19, 8),
    to_signed(22, 8),
    to_signed(17, 8),
    to_signed(3, 8),
    to_signed(-16, 8),
    to_signed(-31, 8),
    to_signed(-40, 8),
    to_signed(-38, 8),
    to_signed(-28, 8),
    to_signed(-12, 8),
    to_signed(7, 8),
    to_signed(24, 8),
    to_signed(39, 8),
    to_signed(48, 8),
    to_signed(48, 8),
    to_signed(37, 8),
    to_signed(23, 8),
    to_signed(13, 8),
    to_signed(8, 8),
    to_signed(5, 8),
    to_signed(7, 8),
    to_signed(14, 8),
    to_signed(22, 8),
    to_signed(26, 8),
    to_signed(22, 8),
    to_signed(11, 8),
    to_signed(-4, 8),
    to_signed(-15, 8),
    to_signed(-13, 8),
    to_signed(2, 8),
    to_signed(21, 8),
    to_signed(39, 8),
    to_signed(50, 8),
    to_signed(51, 8),
    to_signed(43, 8),
    to_signed(31, 8),
    to_signed(21, 8),
    to_signed(18, 8),
    to_signed(24, 8),
    to_signed(39, 8),
    to_signed(58, 8),
    to_signed(71, 8),
    to_signed(73, 8),
    to_signed(59, 8),
    to_signed(24, 8),
    to_signed(-22, 8),
    to_signed(-63, 8),
    to_signed(-83, 8),
    to_signed(-78, 8),
    to_signed(-57, 8),
    to_signed(-31, 8),
    to_signed(-9, 8),
    to_signed(4, 8),
    to_signed(6, 8),
    to_signed(-7, 8),
    to_signed(-30, 8),
    to_signed(-54, 8),
    to_signed(-70, 8),
    to_signed(-74, 8),
    to_signed(-65, 8),
    to_signed(-47, 8),
    to_signed(-26, 8),
    to_signed(-5, 8),
    to_signed(14, 8),
    to_signed(28, 8),
    to_signed(37, 8),
    to_signed(42, 8),
    to_signed(44, 8),
    to_signed(41, 8),
    to_signed(28, 8),
    to_signed(10, 8),
    to_signed(-7, 8),
    to_signed(-19, 8),
    to_signed(-26, 8),
    to_signed(-28, 8),
    to_signed(-22, 8),
    to_signed(-7, 8),
    to_signed(10, 8),
    to_signed(21, 8),
    to_signed(24, 8),
    to_signed(20, 8),
    to_signed(9, 8),
    to_signed(-9, 8),
    to_signed(-29, 8),
    to_signed(-44, 8),
    to_signed(-48, 8),
    to_signed(-40, 8),
    to_signed(-23, 8),
    to_signed(-1, 8),
    to_signed(17, 8),
    to_signed(30, 8),
    to_signed(39, 8),
    to_signed(42, 8),
    to_signed(36, 8),
    to_signed(23, 8),
    to_signed(11, 8),
    to_signed(6, 8),
    to_signed(7, 8),
    to_signed(13, 8),
    to_signed(22, 8),
    to_signed(29, 8),
    to_signed(31, 8),
    to_signed(26, 8),
    to_signed(13, 8),
    to_signed(-4, 8),
    to_signed(-17, 8),
    to_signed(-20, 8),
    to_signed(-10, 8),
    to_signed(8, 8),
    to_signed(26, 8),
    to_signed(38, 8),
    to_signed(38, 8),
    to_signed(29, 8),
    to_signed(15, 8),
    to_signed(3, 8),
    to_signed(-4, 8),
    to_signed(-2, 8),
    to_signed(12, 8),
    to_signed(33, 8),
    to_signed(54, 8),
    to_signed(65, 8),
    to_signed(62, 8),
    to_signed(40, 8),
    to_signed(-1, 8),
    to_signed(-45, 8),
    to_signed(-75, 8),
    to_signed(-83, 8),
    to_signed(-72, 8),
    to_signed(-52, 8),
    to_signed(-30, 8),
    to_signed(-14, 8),
    to_signed(-7, 8),
    to_signed(-12, 8),
    to_signed(-29, 8),
    to_signed(-52, 8),
    to_signed(-70, 8),
    to_signed(-77, 8),
    to_signed(-74, 8),
    to_signed(-64, 8),
    to_signed(-49, 8),
    to_signed(-33, 8),
    to_signed(-18, 8),
    to_signed(-3, 8),
    to_signed(12, 8),
    to_signed(24, 8),
    to_signed(33, 8),
    to_signed(36, 8),
    to_signed(30, 8),
    to_signed(12, 8),
    to_signed(-12, 8),
    to_signed(-29, 8),
    to_signed(-37, 8),
    to_signed(-38, 8),
    to_signed(-32, 8),
    to_signed(-20, 8),
    to_signed(-6, 8),
    to_signed(5, 8),
    to_signed(6, 8),
    to_signed(0, 8),
    to_signed(-11, 8),
    to_signed(-23, 8),
    to_signed(-37, 8),
    to_signed(-47, 8),
    to_signed(-47, 8),
    to_signed(-39, 8),
    to_signed(-26, 8),
    to_signed(-9, 8),
    to_signed(5, 8),
    to_signed(13, 8),
    to_signed(16, 8),
    to_signed(17, 8),
    to_signed(16, 8),
    to_signed(10, 8),
    to_signed(2, 8),
    to_signed(-4, 8),
    to_signed(-4, 8),
    to_signed(2, 8),
    to_signed(13, 8),
    to_signed(24, 8),
    to_signed(28, 8),
    to_signed(22, 8),
    to_signed(9, 8),
    to_signed(-8, 8),
    to_signed(-22, 8),
    to_signed(-26, 8),
    to_signed(-19, 8),
    to_signed(-4, 8),
    to_signed(16, 8),
    to_signed(33, 8),
    to_signed(41, 8),
    to_signed(37, 8),
    to_signed(25, 8),
    to_signed(12, 8),
    to_signed(3, 8),
    to_signed(2, 8),
    to_signed(9, 8),
    to_signed(22, 8),
    to_signed(37, 8),
    to_signed(49, 8),
    to_signed(54, 8),
    to_signed(44, 8),
    to_signed(18, 8),
    to_signed(-19, 8),
    to_signed(-55, 8),
    to_signed(-75, 8),
    to_signed(-75, 8),
    to_signed(-60, 8),
    to_signed(-39, 8),
    to_signed(-19, 8),
    to_signed(-4, 8),
    to_signed(3, 8),
    to_signed(-5, 8),
    to_signed(-25, 8),
    to_signed(-48, 8),
    to_signed(-65, 8),
    to_signed(-70, 8),
    to_signed(-63, 8),
    to_signed(-49, 8),
    to_signed(-30, 8),
    to_signed(-13, 8),
    to_signed(3, 8),
    to_signed(19, 8),
    to_signed(34, 8),
    to_signed(43, 8),
    to_signed(44, 8),
    to_signed(40, 8),
    to_signed(28, 8),
    to_signed(10, 8),
    to_signed(-6, 8),
    to_signed(-12, 8),
    to_signed(-12, 8),
    to_signed(-8, 8),
    to_signed(0, 8),
    to_signed(11, 8),
    to_signed(17, 8),
    to_signed(18, 8),
    to_signed(17, 8),
    to_signed(13, 8),
    to_signed(5, 8),
    to_signed(-7, 8),
    to_signed(-20, 8),
    to_signed(-29, 8),
    to_signed(-31, 8),
    to_signed(-23, 8),
    to_signed(-11, 8),
    to_signed(-1, 8),
    to_signed(6, 8),
    to_signed(11, 8),
    to_signed(13, 8),
    to_signed(14, 8),
    to_signed(12, 8),
    to_signed(8, 8),
    to_signed(4, 8),
    to_signed(3, 8),
    to_signed(5, 8),
    to_signed(10, 8),
    to_signed(17, 8),
    to_signed(21, 8),
    to_signed(19, 8),
    to_signed(11, 8),
    to_signed(-1, 8),
    to_signed(-13, 8),
    to_signed(-21, 8),
    to_signed(-20, 8),
    to_signed(-10, 8),
    to_signed(4, 8),
    to_signed(20, 8),
    to_signed(32, 8),
    to_signed(36, 8),
    to_signed(30, 8),
    to_signed(20, 8),
    to_signed(10, 8),
    to_signed(4, 8),
    to_signed(6, 8),
    to_signed(20, 8),
    to_signed(39, 8),
    to_signed(55, 8),
    to_signed(66, 8),
    to_signed(65, 8),
    to_signed(48, 8),
    to_signed(16, 8),
    to_signed(-21, 8),
    to_signed(-52, 8),
    to_signed(-65, 8),
    to_signed(-56, 8),
    to_signed(-32, 8),
    to_signed(-6, 8),
    to_signed(13, 8),
    to_signed(22, 8),
    to_signed(17, 8),
    to_signed(-2, 8),
    to_signed(-27, 8),
    to_signed(-50, 8),
    to_signed(-63, 8),
    to_signed(-61, 8),
    to_signed(-46, 8),
    to_signed(-24, 8),
    to_signed(-4, 8),
    to_signed(12, 8),
    to_signed(24, 8),
    to_signed(34, 8),
    to_signed(42, 8),
    to_signed(44, 8),
    to_signed(40, 8),
    to_signed(28, 8),
    to_signed(11, 8),
    to_signed(-6, 8),
    to_signed(-16, 8),
    to_signed(-19, 8),
    to_signed(-18, 8),
    to_signed(-17, 8),
    to_signed(-13, 8),
    to_signed(-7, 8),
    to_signed(-4, 8),
    to_signed(-4, 8),
    to_signed(-5, 8),
    to_signed(-8, 8),
    to_signed(-15, 8),
    to_signed(-25, 8),
    to_signed(-33, 8),
    to_signed(-40, 8),
    to_signed(-39, 8),
    to_signed(-30, 8),
    to_signed(-16, 8),
    to_signed(-3, 8),
    to_signed(7, 8),
    to_signed(14, 8),
    to_signed(18, 8),
    to_signed(19, 8),
    to_signed(18, 8),
    to_signed(15, 8),
    to_signed(11, 8),
    to_signed(11, 8),
    to_signed(16, 8),
    to_signed(24, 8),
    to_signed(28, 8),
    to_signed(28, 8),
    to_signed(23, 8),
    to_signed(14, 8),
    to_signed(5, 8),
    to_signed(-1, 8),
    to_signed(-2, 8),
    to_signed(3, 8),
    to_signed(16, 8),
    to_signed(33, 8),
    to_signed(47, 8),
    to_signed(52, 8),
    to_signed(48, 8),
    to_signed(36, 8),
    to_signed(25, 8),
    to_signed(16, 8),
    to_signed(15, 8),
    to_signed(21, 8),
    to_signed(36, 8),
    to_signed(53, 8),
    to_signed(68, 8),
    to_signed(73, 8),
    to_signed(65, 8),
    to_signed(40, 8),
    to_signed(5, 8),
    to_signed(-32, 8),
    to_signed(-60, 8),
    to_signed(-69, 8),
    to_signed(-58, 8),
    to_signed(-37, 8),
    to_signed(-16, 8),
    to_signed(0, 8),
    to_signed(6, 8),
    to_signed(-3, 8),
    to_signed(-24, 8),
    to_signed(-48, 8),
    to_signed(-68, 8),
    to_signed(-82, 8),
    to_signed(-84, 8),
    to_signed(-72, 8),
    to_signed(-54, 8),
    to_signed(-36, 8),
    to_signed(-20, 8),
    to_signed(-6, 8),
    to_signed(5, 8),
    to_signed(13, 8),
    to_signed(18, 8),
    to_signed(20, 8),
    to_signed(15, 8),
    to_signed(5, 8),
    to_signed(-5, 8),
    to_signed(-11, 8),
    to_signed(-14, 8),
    to_signed(-16, 8),
    to_signed(-17, 8),
    to_signed(-16, 8),
    to_signed(-10, 8),
    to_signed(-3, 8),
    to_signed(2, 8),
    to_signed(4, 8),
    to_signed(2, 8),
    to_signed(-7, 8),
    to_signed(-16, 8),
    to_signed(-23, 8),
    to_signed(-26, 8),
    to_signed(-26, 8),
    to_signed(-23, 8),
    to_signed(-15, 8),
    to_signed(-5, 8),
    to_signed(4, 8),
    to_signed(12, 8),
    to_signed(18, 8),
    to_signed(24, 8),
    to_signed(28, 8),
    to_signed(30, 8),
    to_signed(29, 8),
    to_signed(28, 8),
    to_signed(28, 8),
    to_signed(29, 8),
    to_signed(28, 8),
    to_signed(23, 8),
    to_signed(13, 8),
    to_signed(-2, 8),
    to_signed(-15, 8),
    to_signed(-24, 8),
    to_signed(-24, 8),
    to_signed(-15, 8),
    to_signed(2, 8),
    to_signed(19, 8),
    to_signed(30, 8),
    to_signed(33, 8),
    to_signed(26, 8),
    to_signed(11, 8),
    to_signed(-6, 8),
    to_signed(-16, 8),
    to_signed(-15, 8),
    to_signed(-5, 8),
    to_signed(12, 8),
    to_signed(34, 8),
    to_signed(53, 8),
    to_signed(61, 8),
    to_signed(54, 8),
    to_signed(31, 8),
    to_signed(-4, 8),
    to_signed(-43, 8),
    to_signed(-70, 8),
    to_signed(-74, 8),
    to_signed(-62, 8),
    to_signed(-43, 8),
    to_signed(-23, 8),
    to_signed(-5, 8),
    to_signed(2, 8),
    to_signed(-4, 8),
    to_signed(-21, 8),
    to_signed(-38, 8),
    to_signed(-53, 8),
    to_signed(-63, 8),
    to_signed(-62, 8),
    to_signed(-50, 8),
    to_signed(-35, 8),
    to_signed(-22, 8),
    to_signed(-9, 8),
    to_signed(7, 8),
    to_signed(19, 8),
    to_signed(26, 8),
    to_signed(29, 8),
    to_signed(28, 8),
    to_signed(24, 8),
    to_signed(14, 8),
    to_signed(3, 8),
    to_signed(-5, 8),
    to_signed(-11, 8),
    to_signed(-16, 8),
    to_signed(-18, 8),
    to_signed(-15, 8),
    to_signed(-9, 8),
    to_signed(-4, 8),
    to_signed(-1, 8),
    to_signed(1, 8),
    to_signed(-2, 8),
    to_signed(-11, 8),
    to_signed(-22, 8),
    to_signed(-29, 8),
    to_signed(-31, 8),
    to_signed(-29, 8),
    to_signed(-25, 8),
    to_signed(-19, 8),
    to_signed(-11, 8),
    to_signed(-3, 8),
    to_signed(2, 8),
    to_signed(6, 8),
    to_signed(8, 8),
    to_signed(8, 8),
    to_signed(8, 8),
    to_signed(10, 8),
    to_signed(14, 8),
    to_signed(18, 8),
    to_signed(21, 8),
    to_signed(24, 8),
    to_signed(24, 8),
    to_signed(16, 8),
    to_signed(2, 8),
    to_signed(-12, 8),
    to_signed(-21, 8),
    to_signed(-20, 8),
    to_signed(-9, 8),
    to_signed(8, 8),
    to_signed(22, 8),
    to_signed(31, 8),
    to_signed(33, 8),
    to_signed(27, 8),
    to_signed(14, 8),
    to_signed(0, 8),
    to_signed(-9, 8),
    to_signed(-8, 8),
    to_signed(0, 8),
    to_signed(16, 8),
    to_signed(36, 8),
    to_signed(52, 8),
    to_signed(59, 8),
    to_signed(54, 8),
    to_signed(36, 8),
    to_signed(6, 8),
    to_signed(-28, 8),
    to_signed(-50, 8),
    to_signed(-53, 8),
    to_signed(-39, 8),
    to_signed(-18, 8),
    to_signed(1, 8),
    to_signed(13, 8),
    to_signed(14, 8),
    to_signed(3, 8),
    to_signed(-16, 8),
    to_signed(-33, 8),
    to_signed(-47, 8),
    to_signed(-55, 8),
    to_signed(-52, 8),
    to_signed(-40, 8),
    to_signed(-25, 8),
    to_signed(-12, 8),
    to_signed(1, 8),
    to_signed(14, 8),
    to_signed(26, 8),
    to_signed(34, 8),
    to_signed(37, 8),
    to_signed(36, 8),
    to_signed(32, 8),
    to_signed(24, 8),
    to_signed(12, 8),
    to_signed(2, 8),
    to_signed(-5, 8),
    to_signed(-11, 8),
    to_signed(-14, 8),
    to_signed(-11, 8),
    to_signed(-3, 8),
    to_signed(2, 8),
    to_signed(5, 8),
    to_signed(5, 8),
    to_signed(2, 8),
    to_signed(-7, 8),
    to_signed(-19, 8),
    to_signed(-30, 8),
    to_signed(-35, 8),
    to_signed(-34, 8),
    to_signed(-27, 8),
    to_signed(-17, 8),
    to_signed(-8, 8),
    to_signed(1, 8),
    to_signed(7, 8),
    to_signed(11, 8),
    to_signed(13, 8),
    to_signed(12, 8),
    to_signed(10, 8),
    to_signed(8, 8),
    to_signed(10, 8),
    to_signed(12, 8),
    to_signed(12, 8),
    to_signed(13, 8),
    to_signed(13, 8),
    to_signed(11, 8),
    to_signed(5, 8),
    to_signed(-3, 8),
    to_signed(-7, 8),
    to_signed(-3, 8),
    to_signed(11, 8),
    to_signed(29, 8),
    to_signed(44, 8),
    to_signed(53, 8),
    to_signed(54, 8),
    to_signed(46, 8),
    to_signed(34, 8),
    to_signed(23, 8),
    to_signed(18, 8),
    to_signed(20, 8),
    to_signed(29, 8),
    to_signed(44, 8),
    to_signed(60, 8),
    to_signed(73, 8),
    to_signed(75, 8),
    to_signed(64, 8),
    to_signed(37, 8),
    to_signed(2, 8),
    to_signed(-33, 8),
    to_signed(-55, 8),
    to_signed(-57, 8),
    to_signed(-43, 8),
    to_signed(-21, 8),
    to_signed(-1, 8),
    to_signed(13, 8),
    to_signed(17, 8),
    to_signed(8, 8),
    to_signed(-11, 8),
    to_signed(-32, 8),
    to_signed(-48, 8),
    to_signed(-57, 8),
    to_signed(-57, 8),
    to_signed(-46, 8),
    to_signed(-28, 8),
    to_signed(-11, 8),
    to_signed(2, 8),
    to_signed(13, 8),
    to_signed(21, 8),
    to_signed(27, 8),
    to_signed(28, 8),
    to_signed(28, 8),
    to_signed(25, 8),
    to_signed(16, 8),
    to_signed(1, 8),
    to_signed(-9, 8),
    to_signed(-14, 8),
    to_signed(-18, 8),
    to_signed(-23, 8),
    to_signed(-22, 8),
    to_signed(-12, 8),
    to_signed(-3, 8),
    to_signed(3, 8),
    to_signed(5, 8),
    to_signed(2, 8),
    to_signed(-8, 8),
    to_signed(-22, 8),
    to_signed(-32, 8),
    to_signed(-35, 8),
    to_signed(-32, 8),
    to_signed(-23, 8),
    to_signed(-11, 8),
    to_signed(3, 8),
    to_signed(12, 8),
    to_signed(17, 8),
    to_signed(21, 8),
    to_signed(27, 8),
    to_signed(32, 8),
    to_signed(33, 8),
    to_signed(34, 8),
    to_signed(37, 8),
    to_signed(41, 8),
    to_signed(42, 8),
    to_signed(42, 8),
    to_signed(41, 8),
    to_signed(36, 8),
    to_signed(26, 8),
    to_signed(17, 8),
    to_signed(10, 8),
    to_signed(10, 8),
    to_signed(17, 8),
    to_signed(29, 8),
    to_signed(39, 8),
    to_signed(44, 8),
    to_signed(42, 8),
    to_signed(34, 8),
    to_signed(22, 8),
    to_signed(12, 8),
    to_signed(8, 8),
    to_signed(10, 8),
    to_signed(20, 8),
    to_signed(35, 8),
    to_signed(51, 8),
    to_signed(61, 8),
    to_signed(63, 8),
    to_signed(49, 8),
    to_signed(22, 8),
    to_signed(-13, 8),
    to_signed(-44, 8),
    to_signed(-63, 8),
    to_signed(-64, 8),
    to_signed(-52, 8),
    to_signed(-35, 8),
    to_signed(-20, 8),
    to_signed(-7, 8),
    to_signed(-3, 8),
    to_signed(-14, 8),
    to_signed(-35, 8),
    to_signed(-57, 8),
    to_signed(-72, 8),
    to_signed(-76, 8),
    to_signed(-71, 8),
    to_signed(-58, 8),
    to_signed(-41, 8),
    to_signed(-25, 8),
    to_signed(-10, 8),
    to_signed(4, 8),
    to_signed(16, 8),
    to_signed(25, 8),
    to_signed(30, 8),
    to_signed(33, 8),
    to_signed(32, 8),
    to_signed(25, 8),
    to_signed(11, 8),
    to_signed(-1, 8),
    to_signed(-7, 8),
    to_signed(-10, 8),
    to_signed(-14, 8),
    to_signed(-12, 8),
    to_signed(-4, 8),
    to_signed(4, 8),
    to_signed(9, 8),
    to_signed(11, 8),
    to_signed(7, 8),
    to_signed(-4, 8),
    to_signed(-17, 8),
    to_signed(-26, 8),
    to_signed(-29, 8),
    to_signed(-26, 8),
    to_signed(-20, 8),
    to_signed(-11, 8),
    to_signed(-2, 8),
    to_signed(6, 8),
    to_signed(8, 8),
    to_signed(8, 8),
    to_signed(10, 8),
    to_signed(12, 8),
    to_signed(11, 8),
    to_signed(10, 8),
    to_signed(11, 8),
    to_signed(11, 8),
    to_signed(9, 8),
    to_signed(6, 8),
    to_signed(3, 8),
    to_signed(-3, 8),
    to_signed(-10, 8),
    to_signed(-16, 8),
    to_signed(-19, 8),
    to_signed(-18, 8),
    to_signed(-12, 8),
    to_signed(-1, 8),
    to_signed(9, 8),
    to_signed(13, 8),
    to_signed(12, 8),
    to_signed(6, 8),
    to_signed(-5, 8),
    to_signed(-15, 8),
    to_signed(-19, 8),
    to_signed(-15, 8),
    to_signed(-1, 8),
    to_signed(18, 8),
    to_signed(37, 8),
    to_signed(48, 8),
    to_signed(49, 8),
    to_signed(37, 8),
    to_signed(13, 8),
    to_signed(-18, 8),
    to_signed(-46, 8),
    to_signed(-63, 8),
    to_signed(-60, 8),
    to_signed(-43, 8),
    to_signed(-24, 8),
    to_signed(-9, 8),
    to_signed(0, 8),
    to_signed(1, 8),
    to_signed(-10, 8),
    to_signed(-28, 8),
    to_signed(-45, 8),
    to_signed(-56, 8),
    to_signed(-59, 8),
    to_signed(-53, 8),
    to_signed(-44, 8),
    to_signed(-37, 8),
    to_signed(-32, 8),
    to_signed(-23, 8),
    to_signed(-11, 8),
    to_signed(2, 8),
    to_signed(16, 8),
    to_signed(29, 8),
    to_signed(39, 8),
    to_signed(41, 8),
    to_signed(35, 8),
    to_signed(21, 8),
    to_signed(6, 8),
    to_signed(-4, 8),
    to_signed(-10, 8),
    to_signed(-13, 8),
    to_signed(-12, 8),
    to_signed(-7, 8),
    to_signed(-1, 8),
    to_signed(5, 8),
    to_signed(7, 8),
    to_signed(5, 8),
    to_signed(-5, 8),
    to_signed(-18, 8),
    to_signed(-28, 8),
    to_signed(-36, 8),
    to_signed(-37, 8),
    to_signed(-32, 8),
    to_signed(-22, 8),
    to_signed(-10, 8),
    to_signed(2, 8),
    to_signed(12, 8),
    to_signed(18, 8),
    to_signed(22, 8),
    to_signed(25, 8),
    to_signed(27, 8),
    to_signed(27, 8),
    to_signed(30, 8),
    to_signed(31, 8),
    to_signed(28, 8),
    to_signed(24, 8),
    to_signed(21, 8),
    to_signed(18, 8),
    to_signed(14, 8),
    to_signed(12, 8),
    to_signed(10, 8),
    to_signed(7, 8),
    to_signed(9, 8),
    to_signed(17, 8),
    to_signed(27, 8),
    to_signed(31, 8),
    to_signed(28, 8),
    to_signed(22, 8),
    to_signed(13, 8),
    to_signed(4, 8),
    to_signed(-2, 8),
    to_signed(-3, 8),
    to_signed(5, 8),
    to_signed(22, 8),
    to_signed(42, 8),
    to_signed(58, 8),
    to_signed(61, 8),
    to_signed(48, 8),
    to_signed(20, 8),
    to_signed(-13, 8),
    to_signed(-44, 8),
    to_signed(-66, 8),
    to_signed(-71, 8),
    to_signed(-57, 8),
    to_signed(-35, 8),
    to_signed(-18, 8),
    to_signed(-7, 8),
    to_signed(0, 8),
    to_signed(-5, 8),
    to_signed(-20, 8),
    to_signed(-37, 8),
    to_signed(-48, 8),
    to_signed(-52, 8),
    to_signed(-48, 8),
    to_signed(-37, 8),
    to_signed(-25, 8),
    to_signed(-19, 8),
    to_signed(-13, 8),
    to_signed(-5, 8),
    to_signed(7, 8),
    to_signed(20, 8),
    to_signed(30, 8),
    to_signed(38, 8),
    to_signed(40, 8),
    to_signed(30, 8),
    to_signed(13, 8),
    to_signed(-4, 8),
    to_signed(-14, 8),
    to_signed(-18, 8),
    to_signed(-19, 8),
    to_signed(-15, 8),
    to_signed(-6, 8),
    to_signed(1, 8),
    to_signed(5, 8),
    to_signed(7, 8),
    to_signed(5, 8),
    to_signed(-5, 8),
    to_signed(-18, 8),
    to_signed(-27, 8),
    to_signed(-32, 8),
    to_signed(-36, 8),
    to_signed(-33, 8),
    to_signed(-23, 8),
    to_signed(-11, 8),
    to_signed(0, 8),
    to_signed(9, 8),
    to_signed(17, 8),
    to_signed(19, 8),
    to_signed(15, 8),
    to_signed(8, 8),
    to_signed(2, 8),
    to_signed(0, 8),
    to_signed(1, 8),
    to_signed(5, 8),
    to_signed(10, 8),
    to_signed(15, 8),
    to_signed(14, 8),
    to_signed(9, 8),
    to_signed(4, 8),
    to_signed(-2, 8),
    to_signed(-9, 8),
    to_signed(-9, 8),
    to_signed(-1, 8),
    to_signed(10, 8),
    to_signed(16, 8),
    to_signed(18, 8),
    to_signed(17, 8),
    to_signed(10, 8),
    to_signed(0, 8),
    to_signed(-6, 8),
    to_signed(-5, 8),
    to_signed(4, 8),
    to_signed(21, 8),
    to_signed(42, 8),
    to_signed(59, 8),
    to_signed(66, 8),
    to_signed(59, 8),
    to_signed(42, 8),
    to_signed(19, 8),
    to_signed(-6, 8),
    to_signed(-30, 8),
    to_signed(-46, 8),
    to_signed(-47, 8),
    to_signed(-36, 8),
    to_signed(-21, 8),
    to_signed(-6, 8),
    to_signed(4, 8),
    to_signed(6, 8),
    to_signed(-3, 8),
    to_signed(-19, 8),
    to_signed(-36, 8),
    to_signed(-50, 8),
    to_signed(-56, 8),
    to_signed(-51, 8),
    to_signed(-40, 8),
    to_signed(-29, 8),
    to_signed(-19, 8),
    to_signed(-6, 8),
    to_signed(8, 8),
    to_signed(20, 8),
    to_signed(30, 8),
    to_signed(35, 8),
    to_signed(35, 8),
    to_signed(28, 8),
    to_signed(16, 8),
    to_signed(1, 8),
    to_signed(-13, 8),
    to_signed(-24, 8),
    to_signed(-30, 8),
    to_signed(-30, 8),
    to_signed(-25, 8),
    to_signed(-19, 8),
    to_signed(-14, 8),
    to_signed(-10, 8),
    to_signed(-10, 8),
    to_signed(-15, 8),
    to_signed(-22, 8),
    to_signed(-28, 8),
    to_signed(-33, 8),
    to_signed(-37, 8),
    to_signed(-35, 8),
    to_signed(-26, 8),
    to_signed(-16, 8),
    to_signed(-6, 8),
    to_signed(5, 8),
    to_signed(17, 8),
    to_signed(24, 8),
    to_signed(25, 8),
    to_signed(23, 8),
    to_signed(19, 8),
    to_signed(16, 8),
    to_signed(15, 8),
    to_signed(15, 8),
    to_signed(15, 8),
    to_signed(13, 8),
    to_signed(11, 8),
    to_signed(8, 8),
    to_signed(5, 8),
    to_signed(0, 8),
    to_signed(-4, 8),
    to_signed(-2, 8),
    to_signed(8, 8),
    to_signed(20, 8),
    to_signed(29, 8),
    to_signed(34, 8),
    to_signed(33, 8),
    to_signed(24, 8),
    to_signed(11, 8),
    to_signed(-1, 8),
    to_signed(-7, 8),
    to_signed(-4, 8),
    to_signed(10, 8),
    to_signed(32, 8),
    to_signed(51, 8),
    to_signed(60, 8),
    to_signed(58, 8),
    to_signed(46, 8),
    to_signed(24, 8),
    to_signed(-2, 8),
    to_signed(-27, 8),
    to_signed(-48, 8),
    to_signed(-59, 8),
    to_signed(-56, 8),
    to_signed(-43, 8),
    to_signed(-29, 8),
    to_signed(-18, 8),
    to_signed(-12, 8),
    to_signed(-12, 8),
    to_signed(-18, 8),
    to_signed(-29, 8),
    to_signed(-40, 8),
    to_signed(-50, 8),
    to_signed(-55, 8),
    to_signed(-54, 8),
    to_signed(-48, 8),
    to_signed(-39, 8),
    to_signed(-27, 8),
    to_signed(-13, 8),
    to_signed(6, 8),
    to_signed(26, 8),
    to_signed(40, 8),
    to_signed(44, 8),
    to_signed(41, 8),
    to_signed(31, 8),
    to_signed(15, 8),
    to_signed(-2, 8),
    to_signed(-13, 8),
    to_signed(-19, 8),
    to_signed(-21, 8),
    to_signed(-18, 8),
    to_signed(-11, 8),
    to_signed(-5, 8),
    to_signed(-1, 8),
    to_signed(1, 8),
    to_signed(-2, 8),
    to_signed(-9, 8),
    to_signed(-19, 8),
    to_signed(-27, 8),
    to_signed(-32, 8),
    to_signed(-33, 8),
    to_signed(-30, 8),
    to_signed(-23, 8),
    to_signed(-13, 8),
    to_signed(-1, 8),
    to_signed(12, 8),
    to_signed(22, 8),
    to_signed(25, 8),
    to_signed(22, 8),
    to_signed(15, 8),
    to_signed(9, 8),
    to_signed(9, 8),
    to_signed(12, 8),
    to_signed(13, 8),
    to_signed(13, 8),
    to_signed(10, 8),
    to_signed(6, 8),
    to_signed(0, 8),
    to_signed(-8, 8),
    to_signed(-18, 8),
    to_signed(-25, 8),
    to_signed(-22, 8),
    to_signed(-10, 8),
    to_signed(3, 8),
    to_signed(12, 8),
    to_signed(15, 8),
    to_signed(11, 8),
    to_signed(2, 8),
    to_signed(-7, 8),
    to_signed(-11, 8),
    to_signed(-9, 8),
    to_signed(0, 8),
    to_signed(17, 8),
    to_signed(35, 8),
    to_signed(49, 8),
    to_signed(53, 8),
    to_signed(48, 8),
    to_signed(36, 8),
    to_signed(18, 8),
    to_signed(-2, 8),
    to_signed(-20, 8),
    to_signed(-34, 8),
    to_signed(-39, 8),
    to_signed(-36, 8),
    to_signed(-27, 8),
    to_signed(-16, 8),
    to_signed(-8, 8),
    to_signed(-5, 8),
    to_signed(-6, 8),
    to_signed(-12, 8),
    to_signed(-24, 8),
    to_signed(-39, 8),
    to_signed(-50, 8),
    to_signed(-51, 8),
    to_signed(-46, 8),
    to_signed(-36, 8),
    to_signed(-25, 8),
    to_signed(-15, 8),
    to_signed(-4, 8),
    to_signed(11, 8),
    to_signed(26, 8),
    to_signed(35, 8),
    to_signed(36, 8),
    to_signed(33, 8),
    to_signed(25, 8),
    to_signed(13, 8),
    to_signed(-1, 8),
    to_signed(-14, 8),
    to_signed(-23, 8),
    to_signed(-25, 8),
    to_signed(-21, 8),
    to_signed(-13, 8),
    to_signed(-7, 8),
    to_signed(-4, 8),
    to_signed(-3, 8),
    to_signed(-4, 8),
    to_signed(-8, 8),
    to_signed(-16, 8),
    to_signed(-26, 8),
    to_signed(-34, 8),
    to_signed(-38, 8),
    to_signed(-34, 8),
    to_signed(-25, 8),
    to_signed(-12, 8),
    to_signed(-1, 8),
    to_signed(8, 8),
    to_signed(16, 8),
    to_signed(23, 8),
    to_signed(24, 8),
    to_signed(19, 8),
    to_signed(14, 8),
    to_signed(13, 8),
    to_signed(14, 8),
    to_signed(17, 8),
    to_signed(20, 8),
    to_signed(20, 8),
    to_signed(19, 8),
    to_signed(20, 8),
    to_signed(20, 8),
    to_signed(16, 8),
    to_signed(9, 8),
    to_signed(6, 8),
    to_signed(10, 8),
    to_signed(19, 8),
    to_signed(27, 8),
    to_signed(32, 8),
    to_signed(30, 8),
    to_signed(25, 8),
    to_signed(17, 8),
    to_signed(12, 8),
    to_signed(11, 8),
    to_signed(14, 8),
    to_signed(23, 8),
    to_signed(36, 8),
    to_signed(49, 8),
    to_signed(57, 8),
    to_signed(55, 8),
    to_signed(46, 8),
    to_signed(34, 8),
    to_signed(16, 8),
    to_signed(-8, 8),
    to_signed(-30, 8),
    to_signed(-43, 8),
    to_signed(-45, 8),
    to_signed(-37, 8),
    to_signed(-19, 8),
    to_signed(-1, 8),
    to_signed(12, 8),
    to_signed(15, 8),
    to_signed(9, 8),
    to_signed(-6, 8),
    to_signed(-30, 8),
    to_signed(-53, 8),
    to_signed(-65, 8),
    to_signed(-64, 8),
    to_signed(-54, 8),
    to_signed(-39, 8),
    to_signed(-21, 8),
    to_signed(-1, 8),
    to_signed(18, 8),
    to_signed(31, 8),
    to_signed(38, 8),
    to_signed(39, 8),
    to_signed(33, 8),
    to_signed(20, 8),
    to_signed(7, 8),
    to_signed(-5, 8),
    to_signed(-16, 8),
    to_signed(-24, 8),
    to_signed(-22, 8),
    to_signed(-15, 8),
    to_signed(-7, 8),
    to_signed(0, 8),
    to_signed(5, 8),
    to_signed(8, 8),
    to_signed(7, 8),
    to_signed(1, 8),
    to_signed(-7, 8),
    to_signed(-18, 8),
    to_signed(-29, 8),
    to_signed(-37, 8),
    to_signed(-37, 8),
    to_signed(-27, 8),
    to_signed(-12, 8),
    to_signed(4, 8),
    to_signed(17, 8),
    to_signed(25, 8),
    to_signed(27, 8),
    to_signed(25, 8),
    to_signed(23, 8),
    to_signed(20, 8),
    to_signed(14, 8),
    to_signed(11, 8),
    to_signed(13, 8),
    to_signed(18, 8),
    to_signed(21, 8),
    to_signed(23, 8),
    to_signed(26, 8),
    to_signed(25, 8),
    to_signed(18, 8),
    to_signed(10, 8),
    to_signed(5, 8),
    to_signed(4, 8),
    to_signed(8, 8),
    to_signed(16, 8),
    to_signed(23, 8),
    to_signed(25, 8),
    to_signed(23, 8),
    to_signed(19, 8),
    to_signed(13, 8),
    to_signed(5, 8),
    to_signed(1, 8),
    to_signed(6, 8),
    to_signed(22, 8),
    to_signed(39, 8),
    to_signed(47, 8),
    to_signed(46, 8),
    to_signed(42, 8),
    to_signed(34, 8),
    to_signed(21, 8),
    to_signed(3, 8),
    to_signed(-19, 8),
    to_signed(-41, 8),
    to_signed(-53, 8),
    to_signed(-48, 8),
    to_signed(-31, 8),
    to_signed(-12, 8),
    to_signed(4, 8),
    to_signed(16, 8),
    to_signed(16, 8),
    to_signed(3, 8),
    to_signed(-20, 8),
    to_signed(-45, 8),
    to_signed(-62, 8),
    to_signed(-66, 8),
    to_signed(-58, 8),
    to_signed(-45, 8),
    to_signed(-31, 8),
    to_signed(-16, 8),
    to_signed(2, 8),
    to_signed(18, 8),
    to_signed(29, 8),
    to_signed(31, 8),
    to_signed(27, 8),
    to_signed(22, 8),
    to_signed(16, 8),
    to_signed(7, 8),
    to_signed(-6, 8),
    to_signed(-16, 8),
    to_signed(-18, 8),
    to_signed(-12, 8),
    to_signed(-4, 8),
    to_signed(2, 8),
    to_signed(5, 8),
    to_signed(7, 8),
    to_signed(12, 8),
    to_signed(16, 8),
    to_signed(13, 8),
    to_signed(1, 8),
    to_signed(-15, 8),
    to_signed(-30, 8),
    to_signed(-37, 8),
    to_signed(-37, 8),
    to_signed(-31, 8),
    to_signed(-22, 8),
    to_signed(-10, 8),
    to_signed(3, 8),
    to_signed(14, 8),
    to_signed(21, 8),
    to_signed(24, 8),
    to_signed(22, 8),
    to_signed(16, 8),
    to_signed(11, 8),
    to_signed(9, 8),
    to_signed(6, 8),
    to_signed(2, 8),
    to_signed(1, 8),
    to_signed(5, 8),
    to_signed(11, 8),
    to_signed(15, 8),
    to_signed(13, 8),
    to_signed(8, 8),
    to_signed(5, 8),
    to_signed(7, 8),
    to_signed(12, 8),
    to_signed(16, 8),
    to_signed(18, 8),
    to_signed(17, 8),
    to_signed(13, 8),
    to_signed(7, 8),
    to_signed(-2, 8),
    to_signed(-10, 8),
    to_signed(-9, 8),
    to_signed(6, 8),
    to_signed(25, 8),
    to_signed(42, 8),
    to_signed(51, 8),
    to_signed(54, 8),
    to_signed(50, 8),
    to_signed(40, 8),
    to_signed(24, 8),
    to_signed(-4, 8),
    to_signed(-39, 8),
    to_signed(-66, 8),
    to_signed(-72, 8),
    to_signed(-57, 8),
    to_signed(-32, 8),
    to_signed(-6, 8),
    to_signed(13, 8),
    to_signed(19, 8),
    to_signed(11, 8),
    to_signed(-7, 8),
    to_signed(-33, 8),
    to_signed(-59, 8),
    to_signed(-74, 8),
    to_signed(-70, 8),
    to_signed(-52, 8),
    to_signed(-32, 8),
    to_signed(-19, 8),
    to_signed(-9, 8),
    to_signed(2, 8),
    to_signed(13, 8),
    to_signed(22, 8),
    to_signed(27, 8),
    to_signed(30, 8),
    to_signed(26, 8),
    to_signed(16, 8),
    to_signed(4, 8),
    to_signed(-7, 8),
    to_signed(-17, 8),
    to_signed(-22, 8),
    to_signed(-18, 8),
    to_signed(-11, 8),
    to_signed(-5, 8),
    to_signed(1, 8),
    to_signed(11, 8),
    to_signed(20, 8),
    to_signed(22, 8),
    to_signed(16, 8),
    to_signed(4, 8),
    to_signed(-14, 8),
    to_signed(-29, 8),
    to_signed(-37, 8),
    to_signed(-35, 8),
    to_signed(-28, 8),
    to_signed(-20, 8),
    to_signed(-10, 8),
    to_signed(3, 8),
    to_signed(14, 8),
    to_signed(21, 8),
    to_signed(22, 8),
    to_signed(20, 8),
    to_signed(16, 8),
    to_signed(13, 8),
    to_signed(10, 8),
    to_signed(7, 8),
    to_signed(3, 8),
    to_signed(2, 8),
    to_signed(6, 8),
    to_signed(11, 8),
    to_signed(11, 8),
    to_signed(10, 8),
    to_signed(12, 8),
    to_signed(20, 8),
    to_signed(27, 8),
    to_signed(32, 8),
    to_signed(35, 8),
    to_signed(33, 8),
    to_signed(26, 8),
    to_signed(14, 8),
    to_signed(2, 8),
    to_signed(-7, 8),
    to_signed(-10, 8),
    to_signed(-1, 8),
    to_signed(16, 8),
    to_signed(35, 8),
    to_signed(48, 8),
    to_signed(56, 8),
    to_signed(59, 8),
    to_signed(56, 8),
    to_signed(44, 8),
    to_signed(23, 8),
    to_signed(-4, 8),
    to_signed(-32, 8),
    to_signed(-55, 8),
    to_signed(-65, 8),
    to_signed(-58, 8),
    to_signed(-38, 8),
    to_signed(-14, 8),
    to_signed(6, 8),
    to_signed(14, 8),
    to_signed(5, 8),
    to_signed(-19, 8),
    to_signed(-46, 8),
    to_signed(-65, 8),
    to_signed(-71, 8),
    to_signed(-64, 8),
    to_signed(-52, 8),
    to_signed(-40, 8),
    to_signed(-30, 8),
    to_signed(-22, 8),
    to_signed(-15, 8),
    to_signed(-8, 8),
    to_signed(2, 8),
    to_signed(15, 8),
    to_signed(28, 8),
    to_signed(36, 8),
    to_signed(35, 8),
    to_signed(22, 8),
    to_signed(2, 8),
    to_signed(-18, 8),
    to_signed(-31, 8),
    to_signed(-32, 8),
    to_signed(-26, 8),
    to_signed(-14, 8),
    to_signed(1, 8),
    to_signed(17, 8),
    to_signed(28, 8),
    to_signed(31, 8),
    to_signed(24, 8),
    to_signed(9, 8),
    to_signed(-9, 8),
    to_signed(-25, 8),
    to_signed(-33, 8),
    to_signed(-33, 8),
    to_signed(-29, 8),
    to_signed(-21, 8),
    to_signed(-6, 8),
    to_signed(13, 8),
    to_signed(26, 8),
    to_signed(30, 8),
    to_signed(28, 8),
    to_signed(23, 8),
    to_signed(17, 8),
    to_signed(8, 8),
    to_signed(1, 8),
    to_signed(-5, 8),
    to_signed(-7, 8),
    to_signed(-5, 8),
    to_signed(-1, 8),
    to_signed(0, 8),
    to_signed(-5, 8),
    to_signed(-9, 8),
    to_signed(-6, 8),
    to_signed(5, 8),
    to_signed(15, 8),
    to_signed(20, 8),
    to_signed(21, 8),
    to_signed(19, 8),
    to_signed(14, 8),
    to_signed(6, 8),
    to_signed(1, 8),
    to_signed(-1, 8),
    to_signed(2, 8),
    to_signed(11, 8),
    to_signed(25, 8),
    to_signed(39, 8),
    to_signed(48, 8),
    to_signed(51, 8),
    to_signed(52, 8),
    to_signed(50, 8),
    to_signed(43, 8),
    to_signed(30, 8),
    to_signed(13, 8),
    to_signed(-8, 8),
    to_signed(-28, 8),
    to_signed(-40, 8),
    to_signed(-38, 8),
    to_signed(-28, 8),
    to_signed(-16, 8),
    to_signed(-8, 8),
    to_signed(-4, 8),
    to_signed(-6, 8),
    to_signed(-14, 8),
    to_signed(-24, 8),
    to_signed(-33, 8),
    to_signed(-38, 8),
    to_signed(-42, 8),
    to_signed(-40, 8),
    to_signed(-34, 8),
    to_signed(-28, 8),
    to_signed(-23, 8),
    to_signed(-19, 8),
    to_signed(-10, 8),
    to_signed(2, 8),
    to_signed(15, 8),
    to_signed(28, 8),
    to_signed(40, 8),
    to_signed(43, 8),
    to_signed(33, 8),
    to_signed(15, 8),
    to_signed(-3, 8),
    to_signed(-19, 8),
    to_signed(-28, 8),
    to_signed(-29, 8),
    to_signed(-23, 8),
    to_signed(-15, 8),
    to_signed(-4, 8),
    to_signed(8, 8),
    to_signed(16, 8),
    to_signed(13, 8),
    to_signed(-2, 8),
    to_signed(-21, 8),
    to_signed(-33, 8),
    to_signed(-39, 8),
    to_signed(-40, 8),
    to_signed(-36, 8),
    to_signed(-30, 8),
    to_signed(-20, 8),
    to_signed(-9, 8),
    to_signed(7, 8),
    to_signed(23, 8),
    to_signed(32, 8),
    to_signed(33, 8),
    to_signed(29, 8),
    to_signed(22, 8),
    to_signed(13, 8),
    to_signed(6, 8),
    to_signed(3, 8),
    to_signed(3, 8),
    to_signed(3, 8),
    to_signed(3, 8),
    to_signed(7, 8),
    to_signed(10, 8),
    to_signed(11, 8),
    to_signed(10, 8),
    to_signed(11, 8),
    to_signed(11, 8),
    to_signed(10, 8),
    to_signed(8, 8),
    to_signed(7, 8),
    to_signed(7, 8),
    to_signed(7, 8),
    to_signed(11, 8),
    to_signed(18, 8),
    to_signed(25, 8),
    to_signed(33, 8),
    to_signed(42, 8),
    to_signed(50, 8),
    to_signed(54, 8),
    to_signed(53, 8),
    to_signed(53, 8),
    to_signed(52, 8),
    to_signed(48, 8),
    to_signed(37, 8),
    to_signed(19, 8),
    to_signed(-3, 8),
    to_signed(-26, 8),
    to_signed(-42, 8),
    to_signed(-48, 8),
    to_signed(-43, 8),
    to_signed(-35, 8),
    to_signed(-26, 8),
    to_signed(-18, 8),
    to_signed(-12, 8),
    to_signed(-15, 8),
    to_signed(-27, 8),
    to_signed(-43, 8),
    to_signed(-58, 8),
    to_signed(-66, 8),
    to_signed(-64, 8),
    to_signed(-55, 8),
    to_signed(-44, 8),
    to_signed(-32, 8),
    to_signed(-16, 8),
    to_signed(6, 8),
    to_signed(27, 8),
    to_signed(41, 8),
    to_signed(46, 8),
    to_signed(44, 8),
    to_signed(37, 8),
    to_signed(26, 8),
    to_signed(10, 8),
    to_signed(-7, 8),
    to_signed(-21, 8),
    to_signed(-26, 8),
    to_signed(-21, 8),
    to_signed(-8, 8),
    to_signed(5, 8),
    to_signed(14, 8),
    to_signed(19, 8),
    to_signed(20, 8),
    to_signed(14, 8),
    to_signed(1, 8),
    to_signed(-13, 8),
    to_signed(-27, 8),
    to_signed(-36, 8),
    to_signed(-39, 8),
    to_signed(-35, 8),
    to_signed(-26, 8),
    to_signed(-12, 8),
    to_signed(4, 8),
    to_signed(23, 8),
    to_signed(37, 8),
    to_signed(42, 8),
    to_signed(38, 8),
    to_signed(29, 8),
    to_signed(18, 8),
    to_signed(5, 8),
    to_signed(-4, 8),
    to_signed(-5, 8),
    to_signed(0, 8),
    to_signed(6, 8),
    to_signed(10, 8),
    to_signed(10, 8),
    to_signed(5, 8),
    to_signed(-3, 8),
    to_signed(-10, 8),
    to_signed(-12, 8),
    to_signed(-10, 8),
    to_signed(-4, 8),
    to_signed(1, 8),
    to_signed(5, 8),
    to_signed(4, 8),
    to_signed(0, 8),
    to_signed(-2, 8),
    to_signed(2, 8),
    to_signed(7, 8),
    to_signed(11, 8),
    to_signed(18, 8),
    to_signed(27, 8),
    to_signed(37, 8),
    to_signed(44, 8),
    to_signed(51, 8),
    to_signed(60, 8),
    to_signed(64, 8),
    to_signed(56, 8),
    to_signed(32, 8),
    to_signed(-3, 8),
    to_signed(-38, 8),
    to_signed(-61, 8),
    to_signed(-66, 8),
    to_signed(-54, 8),
    to_signed(-33, 8),
    to_signed(-12, 8),
    to_signed(5, 8),
    to_signed(12, 8),
    to_signed(4, 8),
    to_signed(-20, 8),
    to_signed(-51, 8),
    to_signed(-74, 8),
    to_signed(-84, 8),
    to_signed(-81, 8),
    to_signed(-67, 8),
    to_signed(-46, 8),
    to_signed(-23, 8),
    to_signed(-1, 8),
    to_signed(22, 8),
    to_signed(44, 8),
    to_signed(57, 8),
    to_signed(56, 8),
    to_signed(45, 8),
    to_signed(28, 8),
    to_signed(9, 8),
    to_signed(-8, 8),
    to_signed(-18, 8),
    to_signed(-18, 8),
    to_signed(-14, 8),
    to_signed(-8, 8),
    to_signed(-1, 8),
    to_signed(7, 8),
    to_signed(11, 8),
    to_signed(10, 8),
    to_signed(4, 8),
    to_signed(-5, 8),
    to_signed(-20, 8),
    to_signed(-37, 8),
    to_signed(-47, 8),
    to_signed(-49, 8),
    to_signed(-46, 8),
    to_signed(-37, 8),
    to_signed(-21, 8),
    to_signed(-2, 8),
    to_signed(11, 8),
    to_signed(17, 8),
    to_signed(21, 8),
    to_signed(22, 8),
    to_signed(20, 8),
    to_signed(17, 8),
    to_signed(16, 8),
    to_signed(18, 8),
    to_signed(19, 8),
    to_signed(19, 8),
    to_signed(18, 8),
    to_signed(14, 8),
    to_signed(7, 8),
    to_signed(0, 8),
    to_signed(-4, 8),
    to_signed(-7, 8),
    to_signed(-10, 8),
    to_signed(-10, 8),
    to_signed(-3, 8),
    to_signed(6, 8),
    to_signed(13, 8),
    to_signed(14, 8),
    to_signed(11, 8),
    to_signed(5, 8),
    to_signed(-5, 8),
    to_signed(-12, 8),
    to_signed(-12, 8),
    to_signed(-5, 8),
    to_signed(6, 8),
    to_signed(22, 8),
    to_signed(41, 8),
    to_signed(57, 8),
    to_signed(66, 8),
    to_signed(64, 8),
    to_signed(55, 8),
    to_signed(39, 8),
    to_signed(17, 8),
    to_signed(-7, 8),
    to_signed(-31, 8),
    to_signed(-47, 8),
    to_signed(-52, 8),
    to_signed(-44, 8),
    to_signed(-27, 8),
    to_signed(-11, 8),
    to_signed(-2, 8),
    to_signed(-4, 8),
    to_signed(-16, 8),
    to_signed(-37, 8),
    to_signed(-63, 8),
    to_signed(-84, 8),
    to_signed(-95, 8),
    to_signed(-93, 8),
    to_signed(-80, 8),
    to_signed(-58, 8),
    to_signed(-33, 8),
    to_signed(-11, 8),
    to_signed(3, 8),
    to_signed(12, 8),
    to_signed(17, 8),
    to_signed(20, 8),
    to_signed(20, 8),
    to_signed(16, 8),
    to_signed(7, 8),
    to_signed(-4, 8),
    to_signed(-13, 8),
    to_signed(-17, 8),
    to_signed(-17, 8),
    to_signed(-16, 8),
    to_signed(-12, 8),
    to_signed(-3, 8),
    to_signed(5, 8),
    to_signed(7, 8),
    to_signed(2, 8),
    to_signed(-6, 8),
    to_signed(-14, 8),
    to_signed(-22, 8),
    to_signed(-32, 8),
    to_signed(-42, 8),
    to_signed(-49, 8),
    to_signed(-48, 8),
    to_signed(-38, 8),
    to_signed(-22, 8),
    to_signed(-5, 8),
    to_signed(10, 8),
    to_signed(22, 8),
    to_signed(31, 8),
    to_signed(35, 8),
    to_signed(31, 8),
    to_signed(23, 8),
    to_signed(15, 8),
    to_signed(9, 8),
    to_signed(5, 8),
    to_signed(4, 8),
    to_signed(4, 8),
    to_signed(4, 8),
    to_signed(2, 8),
    to_signed(-3, 8),
    to_signed(-8, 8),
    to_signed(-9, 8),
    to_signed(-7, 8),
    to_signed(0, 8),
    to_signed(8, 8),
    to_signed(12, 8),
    to_signed(9, 8),
    to_signed(0, 8),
    to_signed(-11, 8),
    to_signed(-20, 8),
    to_signed(-25, 8),
    to_signed(-21, 8),
    to_signed(-9, 8),
    to_signed(9, 8),
    to_signed(29, 8),
    to_signed(47, 8),
    to_signed(56, 8),
    to_signed(56, 8),
    to_signed(48, 8),
    to_signed(40, 8),
    to_signed(34, 8),
    to_signed(30, 8),
    to_signed(25, 8),
    to_signed(15, 8),
    to_signed(-2, 8),
    to_signed(-24, 8),
    to_signed(-40, 8),
    to_signed(-43, 8),
    to_signed(-34, 8),
    to_signed(-22, 8),
    to_signed(-12, 8),
    to_signed(-8, 8),
    to_signed(-12, 8),
    to_signed(-24, 8),
    to_signed(-43, 8),
    to_signed(-62, 8),
    to_signed(-77, 8),
    to_signed(-79, 8),
    to_signed(-67, 8),
    to_signed(-47, 8),
    to_signed(-29, 8),
    to_signed(-15, 8),
    to_signed(-3, 8),
    to_signed(9, 8),
    to_signed(18, 8),
    to_signed(24, 8),
    to_signed(29, 8),
    to_signed(33, 8),
    to_signed(32, 8),
    to_signed(24, 8),
    to_signed(11, 8),
    to_signed(-3, 8),
    to_signed(-12, 8),
    to_signed(-14, 8),
    to_signed(-7, 8),
    to_signed(3, 8),
    to_signed(13, 8),
    to_signed(21, 8),
    to_signed(23, 8),
    to_signed(20, 8),
    to_signed(9, 8),
    to_signed(-7, 8),
    to_signed(-22, 8),
    to_signed(-34, 8),
    to_signed(-40, 8),
    to_signed(-40, 8),
    to_signed(-33, 8),
    to_signed(-20, 8),
    to_signed(-6, 8),
    to_signed(9, 8),
    to_signed(22, 8),
    to_signed(35, 8),
    to_signed(43, 8),
    to_signed(43, 8),
    to_signed(33, 8),
    to_signed(20, 8),
    to_signed(9, 8),
    to_signed(2, 8),
    to_signed(0, 8),
    to_signed(2, 8),
    to_signed(6, 8),
    to_signed(10, 8),
    to_signed(13, 8),
    to_signed(15, 8),
    to_signed(13, 8),
    to_signed(7, 8),
    to_signed(1, 8),
    to_signed(-2, 8),
    to_signed(-1, 8),
    to_signed(1, 8),
    to_signed(1, 8),
    to_signed(-2, 8),
    to_signed(-6, 8),
    to_signed(-9, 8),
    to_signed(-5, 8),
    to_signed(4, 8),
    to_signed(15, 8),
    to_signed(24, 8),
    to_signed(32, 8),
    to_signed(40, 8),
    to_signed(47, 8),
    to_signed(52, 8),
    to_signed(56, 8),
    to_signed(58, 8),
    to_signed(55, 8),
    to_signed(44, 8),
    to_signed(27, 8),
    to_signed(7, 8),
    to_signed(-14, 8),
    to_signed(-32, 8),
    to_signed(-40, 8),
    to_signed(-36, 8),
    to_signed(-23, 8),
    to_signed(-8, 8),
    to_signed(5, 8),
    to_signed(10, 8),
    to_signed(2, 8),
    to_signed(-16, 8),
    to_signed(-38, 8),
    to_signed(-57, 8),
    to_signed(-69, 8),
    to_signed(-71, 8),
    to_signed(-61, 8),
    to_signed(-45, 8),
    to_signed(-29, 8),
    to_signed(-16, 8),
    to_signed(-2, 8),
    to_signed(9, 8),
    to_signed(17, 8),
    to_signed(20, 8),
    to_signed(22, 8),
    to_signed(21, 8),
    to_signed(16, 8),
    to_signed(5, 8),
    to_signed(-6, 8),
    to_signed(-15, 8),
    to_signed(-20, 8),
    to_signed(-18, 8),
    to_signed(-8, 8),
    to_signed(5, 8),
    to_signed(16, 8),
    to_signed(24, 8),
    to_signed(25, 8),
    to_signed(19, 8),
    to_signed(6, 8),
    to_signed(-9, 8),
    to_signed(-21, 8),
    to_signed(-29, 8),
    to_signed(-32, 8),
    to_signed(-30, 8),
    to_signed(-20, 8),
    to_signed(-7, 8),
    to_signed(6, 8),
    to_signed(20, 8),
    to_signed(32, 8),
    to_signed(39, 8),
    to_signed(40, 8),
    to_signed(36, 8),
    to_signed(30, 8),
    to_signed(25, 8),
    to_signed(22, 8),
    to_signed(20, 8),
    to_signed(17, 8),
    to_signed(13, 8),
    to_signed(10, 8),
    to_signed(10, 8),
    to_signed(12, 8),
    to_signed(11, 8),
    to_signed(9, 8),
    to_signed(8, 8),
    to_signed(9, 8),
    to_signed(10, 8),
    to_signed(9, 8),
    to_signed(4, 8),
    to_signed(-2, 8),
    to_signed(-8, 8),
    to_signed(-10, 8),
    to_signed(-7, 8),
    to_signed(0, 8),
    to_signed(11, 8),
    to_signed(26, 8),
    to_signed(41, 8),
    to_signed(51, 8),
    to_signed(55, 8),
    to_signed(53, 8),
    to_signed(48, 8),
    to_signed(43, 8),
    to_signed(40, 8),
    to_signed(39, 8),
    to_signed(38, 8),
    to_signed(30, 8),
    to_signed(15, 8),
    to_signed(-7, 8),
    to_signed(-32, 8),
    to_signed(-50, 8),
    to_signed(-53, 8),
    to_signed(-41, 8),
    to_signed(-22, 8),
    to_signed(-5, 8),
    to_signed(4, 8),
    to_signed(0, 8),
    to_signed(-16, 8),
    to_signed(-40, 8),
    to_signed(-63, 8),
    to_signed(-76, 8),
    to_signed(-74, 8),
    to_signed(-59, 8),
    to_signed(-36, 8),
    to_signed(-16, 8),
    to_signed(-3, 8),
    to_signed(5, 8),
    to_signed(14, 8),
    to_signed(24, 8),
    to_signed(32, 8),
    to_signed(36, 8),
    to_signed(38, 8),
    to_signed(37, 8),
    to_signed(29, 8),
    to_signed(16, 8),
    to_signed(3, 8),
    to_signed(-5, 8),
    to_signed(-7, 8),
    to_signed(-2, 8),
    to_signed(6, 8),
    to_signed(15, 8),
    to_signed(21, 8),
    to_signed(26, 8),
    to_signed(29, 8),
    to_signed(27, 8),
    to_signed(15, 8),
    to_signed(-3, 8),
    to_signed(-18, 8),
    to_signed(-27, 8),
    to_signed(-32, 8),
    to_signed(-32, 8),
    to_signed(-24, 8),
    to_signed(-10, 8),
    to_signed(7, 8),
    to_signed(25, 8),
    to_signed(41, 8),
    to_signed(47, 8),
    to_signed(42, 8),
    to_signed(33, 8),
    to_signed(24, 8),
    to_signed(15, 8),
    to_signed(7, 8),
    to_signed(2, 8),
    to_signed(3, 8),
    to_signed(9, 8),
    to_signed(16, 8),
    to_signed(20, 8),
    to_signed(18, 8),
    to_signed(9, 8),
    to_signed(-4, 8),
    to_signed(-13, 8),
    to_signed(-14, 8),
    to_signed(-11, 8),
    to_signed(-6, 8),
    to_signed(-2, 8),
    to_signed(1, 8),
    to_signed(0, 8),
    to_signed(-4, 8),
    to_signed(-7, 8),
    to_signed(-6, 8),
    to_signed(3, 8),
    to_signed(18, 8),
    to_signed(34, 8),
    to_signed(46, 8),
    to_signed(50, 8),
    to_signed(48, 8),
    to_signed(44, 8),
    to_signed(43, 8),
    to_signed(43, 8),
    to_signed(44, 8),
    to_signed(43, 8),
    to_signed(38, 8),
    to_signed(27, 8),
    to_signed(7, 8),
    to_signed(-18, 8),
    to_signed(-40, 8),
    to_signed(-51, 8),
    to_signed(-46, 8),
    to_signed(-28, 8),
    to_signed(-8, 8),
    to_signed(2, 8),
    to_signed(-2, 8),
    to_signed(-17, 8),
    to_signed(-38, 8),
    to_signed(-60, 8),
    to_signed(-78, 8),
    to_signed(-84, 8),
    to_signed(-77, 8),
    to_signed(-55, 8),
    to_signed(-25, 8),
    to_signed(2, 8),
    to_signed(19, 8),
    to_signed(25, 8),
    to_signed(25, 8),
    to_signed(23, 8),
    to_signed(19, 8),
    to_signed(14, 8),
    to_signed(10, 8),
    to_signed(3, 8),
    to_signed(-6, 8),
    to_signed(-15, 8),
    to_signed(-21, 8),
    to_signed(-22, 8),
    to_signed(-16, 8),
    to_signed(-4, 8),
    to_signed(11, 8),
    to_signed(20, 8),
    to_signed(20, 8),
    to_signed(14, 8),
    to_signed(5, 8),
    to_signed(-8, 8),
    to_signed(-20, 8),
    to_signed(-30, 8),
    to_signed(-36, 8),
    to_signed(-37, 8),
    to_signed(-29, 8),
    to_signed(-13, 8),
    to_signed(3, 8),
    to_signed(14, 8),
    to_signed(22, 8),
    to_signed(28, 8),
    to_signed(29, 8),
    to_signed(21, 8),
    to_signed(10, 8),
    to_signed(1, 8),
    to_signed(-4, 8),
    to_signed(-1, 8),
    to_signed(8, 8),
    to_signed(18, 8),
    to_signed(22, 8),
    to_signed(22, 8),
    to_signed(20, 8),
    to_signed(13, 8),
    to_signed(-1, 8),
    to_signed(-14, 8),
    to_signed(-18, 8),
    to_signed(-13, 8),
    to_signed(-3, 8),
    to_signed(5, 8),
    to_signed(10, 8),
    to_signed(9, 8),
    to_signed(-1, 8),
    to_signed(-12, 8),
    to_signed(-20, 8),
    to_signed(-22, 8),
    to_signed(-17, 8),
    to_signed(-4, 8),
    to_signed(15, 8),
    to_signed(30, 8),
    to_signed(37, 8),
    to_signed(37, 8),
    to_signed(33, 8),
    to_signed(24, 8),
    to_signed(17, 8),
    to_signed(15, 8),
    to_signed(20, 8),
    to_signed(24, 8),
    to_signed(22, 8),
    to_signed(10, 8),
    to_signed(-12, 8),
    to_signed(-38, 8),
    to_signed(-55, 8),
    to_signed(-55, 8),
    to_signed(-41, 8),
    to_signed(-23, 8),
    to_signed(-10, 8),
    to_signed(-8, 8),
    to_signed(-17, 8),
    to_signed(-37, 8),
    to_signed(-61, 8),
    to_signed(-79, 8),
    to_signed(-85, 8),
    to_signed(-77, 8),
    to_signed(-57, 8),
    to_signed(-31, 8),
    to_signed(-11, 8),
    to_signed(0, 8),
    to_signed(3, 8),
    to_signed(3, 8),
    to_signed(1, 8),
    to_signed(1, 8),
    to_signed(4, 8),
    to_signed(11, 8),
    to_signed(17, 8),
    to_signed(15, 8),
    to_signed(6, 8),
    to_signed(-5, 8),
    to_signed(-14, 8),
    to_signed(-17, 8),
    to_signed(-11, 8),
    to_signed(1, 8),
    to_signed(12, 8),
    to_signed(17, 8),
    to_signed(18, 8),
    to_signed(15, 8),
    to_signed(7, 8),
    to_signed(-7, 8),
    to_signed(-20, 8),
    to_signed(-28, 8),
    to_signed(-31, 8),
    to_signed(-27, 8),
    to_signed(-19, 8),
    to_signed(-9, 8),
    to_signed(-3, 8),
    to_signed(3, 8),
    to_signed(14, 8),
    to_signed(24, 8),
    to_signed(25, 8),
    to_signed(17, 8),
    to_signed(7, 8),
    to_signed(-1, 8),
    to_signed(-8, 8),
    to_signed(-12, 8),
    to_signed(-9, 8),
    to_signed(-4, 8),
    to_signed(2, 8),
    to_signed(7, 8),
    to_signed(9, 8),
    to_signed(5, 8),
    to_signed(-6, 8),
    to_signed(-17, 8),
    to_signed(-21, 8),
    to_signed(-20, 8),
    to_signed(-16, 8),
    to_signed(-10, 8),
    to_signed(-3, 8),
    to_signed(-2, 8),
    to_signed(-8, 8),
    to_signed(-13, 8),
    to_signed(-14, 8),
    to_signed(-13, 8),
    to_signed(-11, 8),
    to_signed(-4, 8),
    to_signed(8, 8),
    to_signed(18, 8),
    to_signed(23, 8),
    to_signed(25, 8),
    to_signed(26, 8),
    to_signed(27, 8),
    to_signed(26, 8),
    to_signed(26, 8),
    to_signed(27, 8),
    to_signed(28, 8),
    to_signed(29, 8),
    to_signed(25, 8),
    to_signed(13, 8),
    to_signed(-9, 8),
    to_signed(-32, 8),
    to_signed(-42, 8),
    to_signed(-37, 8),
    to_signed(-25, 8),
    to_signed(-13, 8),
    to_signed(-4, 8),
    to_signed(0, 8),
    to_signed(-6, 8),
    to_signed(-24, 8),
    to_signed(-47, 8),
    to_signed(-66, 8),
    to_signed(-74, 8),
    to_signed(-66, 8),
    to_signed(-45, 8),
    to_signed(-18, 8),
    to_signed(0, 8),
    to_signed(6, 8),
    to_signed(6, 8),
    to_signed(3, 8),
    to_signed(-1, 8),
    to_signed(-4, 8),
    to_signed(-4, 8),
    to_signed(-1, 8),
    to_signed(1, 8),
    to_signed(1, 8),
    to_signed(-3, 8),
    to_signed(-12, 8),
    to_signed(-22, 8),
    to_signed(-27, 8),
    to_signed(-23, 8),
    to_signed(-13, 8),
    to_signed(-3, 8),
    to_signed(4, 8),
    to_signed(10, 8),
    to_signed(10, 8),
    to_signed(3, 8),
    to_signed(-7, 8),
    to_signed(-15, 8),
    to_signed(-20, 8),
    to_signed(-23, 8),
    to_signed(-21, 8),
    to_signed(-14, 8),
    to_signed(-1, 8),
    to_signed(13, 8),
    to_signed(27, 8),
    to_signed(38, 8),
    to_signed(41, 8),
    to_signed(37, 8),
    to_signed(27, 8),
    to_signed(14, 8),
    to_signed(4, 8),
    to_signed(1, 8),
    to_signed(7, 8),
    to_signed(17, 8),
    to_signed(25, 8),
    to_signed(28, 8),
    to_signed(26, 8),
    to_signed(19, 8),
    to_signed(8, 8),
    to_signed(-5, 8),
    to_signed(-13, 8),
    to_signed(-12, 8),
    to_signed(-1, 8),
    to_signed(10, 8),
    to_signed(16, 8),
    to_signed(12, 8),
    to_signed(0, 8),
    to_signed(-15, 8),
    to_signed(-30, 8),
    to_signed(-37, 8),
    to_signed(-33, 8),
    to_signed(-20, 8),
    to_signed(-3, 8),
    to_signed(11, 8),
    to_signed(19, 8),
    to_signed(19, 8),
    to_signed(14, 8),
    to_signed(6, 8),
    to_signed(2, 8),
    to_signed(3, 8),
    to_signed(10, 8),
    to_signed(19, 8),
    to_signed(25, 8),
    to_signed(22, 8),
    to_signed(12, 8),
    to_signed(-1, 8),
    to_signed(-16, 8),
    to_signed(-31, 8),
    to_signed(-40, 8),
    to_signed(-36, 8),
    to_signed(-21, 8),
    to_signed(-6, 8),
    to_signed(-2, 8),
    to_signed(-10, 8),
    to_signed(-24, 8),
    to_signed(-38, 8),
    to_signed(-51, 8),
    to_signed(-57, 8),
    to_signed(-56, 8),
    to_signed(-46, 8),
    to_signed(-31, 8),
    to_signed(-14, 8),
    to_signed(-1, 8),
    to_signed(3, 8),
    to_signed(3, 8),
    to_signed(4, 8),
    to_signed(10, 8),
    to_signed(18, 8),
    to_signed(25, 8),
    to_signed(30, 8),
    to_signed(29, 8),
    to_signed(22, 8),
    to_signed(11, 8),
    to_signed(2, 8),
    to_signed(-3, 8),
    to_signed(-3, 8),
    to_signed(1, 8),
    to_signed(10, 8),
    to_signed(17, 8),
    to_signed(16, 8),
    to_signed(7, 8),
    to_signed(-4, 8),
    to_signed(-13, 8),
    to_signed(-19, 8),
    to_signed(-22, 8),
    to_signed(-23, 8),
    to_signed(-22, 8),
    to_signed(-19, 8),
    to_signed(-15, 8),
    to_signed(-10, 8),
    to_signed(-5, 8),
    to_signed(3, 8),
    to_signed(12, 8),
    to_signed(18, 8),
    to_signed(19, 8),
    to_signed(17, 8),
    to_signed(12, 8),
    to_signed(6, 8),
    to_signed(-3, 8),
    to_signed(-7, 8),
    to_signed(-3, 8),
    to_signed(5, 8),
    to_signed(12, 8),
    to_signed(13, 8),
    to_signed(8, 8),
    to_signed(-1, 8),
    to_signed(-11, 8),
    to_signed(-18, 8),
    to_signed(-20, 8),
    to_signed(-18, 8),
    to_signed(-11, 8),
    to_signed(-4, 8),
    to_signed(-4, 8),
    to_signed(-10, 8),
    to_signed(-17, 8),
    to_signed(-20, 8),
    to_signed(-19, 8),
    to_signed(-15, 8),
    to_signed(-6, 8),
    to_signed(8, 8),
    to_signed(21, 8),
    to_signed(28, 8),
    to_signed(28, 8),
    to_signed(25, 8),
    to_signed(21, 8),
    to_signed(20, 8),
    to_signed(25, 8),
    to_signed(35, 8),
    to_signed(44, 8),
    to_signed(50, 8),
    to_signed(52, 8),
    to_signed(49, 8),
    to_signed(40, 8),
    to_signed(28, 8),
    to_signed(15, 8),
    to_signed(1, 8),
    to_signed(-12, 8),
    to_signed(-19, 8),
    to_signed(-17, 8),
    to_signed(-10, 8),
    to_signed(-7, 8),
    to_signed(-9, 8),
    to_signed(-12, 8),
    to_signed(-19, 8),
    to_signed(-29, 8),
    to_signed(-39, 8),
    to_signed(-45, 8),
    to_signed(-44, 8),
    to_signed(-36, 8),
    to_signed(-22, 8),
    to_signed(-6, 8),
    to_signed(4, 8),
    to_signed(7, 8),
    to_signed(6, 8),
    to_signed(6, 8),
    to_signed(6, 8),
    to_signed(8, 8),
    to_signed(15, 8),
    to_signed(23, 8),
    to_signed(25, 8),
    to_signed(18, 8),
    to_signed(8, 8),
    to_signed(0, 8),
    to_signed(-7, 8),
    to_signed(-10, 8),
    to_signed(-7, 8),
    to_signed(1, 8),
    to_signed(7, 8),
    to_signed(10, 8),
    to_signed(9, 8),
    to_signed(4, 8),
    to_signed(-7, 8),
    to_signed(-18, 8),
    to_signed(-20, 8),
    to_signed(-17, 8),
    to_signed(-11, 8),
    to_signed(-5, 8),
    to_signed(4, 8),
    to_signed(13, 8),
    to_signed(19, 8),
    to_signed(23, 8),
    to_signed(27, 8),
    to_signed(30, 8),
    to_signed(28, 8),
    to_signed(23, 8),
    to_signed(17, 8),
    to_signed(9, 8),
    to_signed(1, 8),
    to_signed(-1, 8),
    to_signed(6, 8),
    to_signed(15, 8),
    to_signed(18, 8),
    to_signed(16, 8),
    to_signed(11, 8),
    to_signed(5, 8),
    to_signed(-1, 8),
    to_signed(-5, 8),
    to_signed(-3, 8),
    to_signed(-1, 8),
    to_signed(-1, 8),
    to_signed(-2, 8),
    to_signed(-6, 8),
    to_signed(-12, 8),
    to_signed(-17, 8),
    to_signed(-15, 8),
    to_signed(-7, 8),
    to_signed(3, 8),
    to_signed(13, 8),
    to_signed(24, 8),
    to_signed(30, 8),
    to_signed(29, 8),
    to_signed(22, 8),
    to_signed(15, 8),
    to_signed(12, 8),
    to_signed(13, 8),
    to_signed(19, 8),
    to_signed(27, 8),
    to_signed(32, 8),
    to_signed(33, 8),
    to_signed(30, 8),
    to_signed(27, 8),
    to_signed(24, 8),
    to_signed(19, 8),
    to_signed(10, 8),
    to_signed(-3, 8),
    to_signed(-19, 8),
    to_signed(-35, 8),
    to_signed(-44, 8),
    to_signed(-45, 8),
    to_signed(-41, 8),
    to_signed(-37, 8),
    to_signed(-32, 8),
    to_signed(-28, 8),
    to_signed(-27, 8),
    to_signed(-32, 8),
    to_signed(-38, 8),
    to_signed(-42, 8),
    to_signed(-42, 8),
    to_signed(-37, 8),
    to_signed(-24, 8),
    to_signed(-10, 8),
    to_signed(1, 8),
    to_signed(8, 8),
    to_signed(12, 8),
    to_signed(14, 8),
    to_signed(13, 8),
    to_signed(12, 8),
    to_signed(12, 8),
    to_signed(15, 8),
    to_signed(16, 8),
    to_signed(14, 8),
    to_signed(10, 8),
    to_signed(5, 8),
    to_signed(-1, 8),
    to_signed(-4, 8),
    to_signed(-2, 8),
    to_signed(3, 8),
    to_signed(6, 8),
    to_signed(7, 8),
    to_signed(5, 8),
    to_signed(3, 8),
    to_signed(2, 8),
    to_signed(1, 8),
    to_signed(-1, 8),
    to_signed(-3, 8),
    to_signed(-5, 8),
    to_signed(-5, 8),
    to_signed(-1, 8),
    to_signed(2, 8),
    to_signed(3, 8),
    to_signed(6, 8),
    to_signed(10, 8),
    to_signed(14, 8),
    to_signed(13, 8),
    to_signed(6, 8),
    to_signed(-3, 8),
    to_signed(-8, 8),
    to_signed(-11, 8),
    to_signed(-11, 8),
    to_signed(-8, 8),
    to_signed(-3, 8),
    to_signed(2, 8),
    to_signed(1, 8),
    to_signed(-6, 8),
    to_signed(-17, 8),
    to_signed(-27, 8),
    to_signed(-30, 8),
    to_signed(-26, 8),
    to_signed(-17, 8),
    to_signed(-8, 8),
    to_signed(-4, 8),
    to_signed(-3, 8),
    to_signed(-4, 8),
    to_signed(-8, 8),
    to_signed(-12, 8),
    to_signed(-13, 8),
    to_signed(-10, 8),
    to_signed(-2, 8),
    to_signed(10, 8),
    to_signed(21, 8),
    to_signed(28, 8),
    to_signed(30, 8),
    to_signed(31, 8),
    to_signed(34, 8),
    to_signed(35, 8),
    to_signed(33, 8),
    to_signed(29, 8),
    to_signed(26, 8),
    to_signed(25, 8),
    to_signed(26, 8),
    to_signed(27, 8),
    to_signed(29, 8),
    to_signed(29, 8),
    to_signed(24, 8),
    to_signed(14, 8),
    to_signed(2, 8),
    to_signed(-11, 8),
    to_signed(-22, 8),
    to_signed(-26, 8),
    to_signed(-22, 8),
    to_signed(-15, 8),
    to_signed(-6, 8),
    to_signed(0, 8),
    to_signed(-2, 8),
    to_signed(-13, 8),
    to_signed(-27, 8),
    to_signed(-35, 8),
    to_signed(-35, 8),
    to_signed(-29, 8),
    to_signed(-18, 8),
    to_signed(-5, 8),
    to_signed(4, 8),
    to_signed(4, 8),
    to_signed(-3, 8),
    to_signed(-11, 8),
    to_signed(-16, 8),
    to_signed(-16, 8),
    to_signed(-11, 8),
    to_signed(-2, 8),
    to_signed(3, 8),
    to_signed(4, 8),
    to_signed(1, 8),
    to_signed(-5, 8),
    to_signed(-11, 8),
    to_signed(-13, 8),
    to_signed(-10, 8),
    to_signed(-3, 8),
    to_signed(2, 8),
    to_signed(6, 8),
    to_signed(8, 8),
    to_signed(6, 8),
    to_signed(1, 8),
    to_signed(-4, 8),
    to_signed(-5, 8),
    to_signed(-1, 8),
    to_signed(5, 8),
    to_signed(7, 8),
    to_signed(7, 8),
    to_signed(5, 8),
    to_signed(4, 8),
    to_signed(4, 8),
    to_signed(3, 8),
    to_signed(1, 8),
    to_signed(0, 8),
    to_signed(1, 8),
    to_signed(5, 8),
    to_signed(9, 8),
    to_signed(14, 8),
    to_signed(19, 8),
    to_signed(24, 8),
    to_signed(26, 8),
    to_signed(22, 8),
    to_signed(13, 8),
    to_signed(2, 8),
    to_signed(-6, 8),
    to_signed(-9, 8),
    to_signed(-9, 8),
    to_signed(-5, 8),
    to_signed(1, 8),
    to_signed(6, 8),
    to_signed(8, 8),
    to_signed(5, 8),
    to_signed(-1, 8),
    to_signed(-8, 8),
    to_signed(-14, 8),
    to_signed(-16, 8),
    to_signed(-14, 8),
    to_signed(-10, 8),
    to_signed(-7, 8),
    to_signed(-3, 8),
    to_signed(2, 8),
    to_signed(7, 8),
    to_signed(12, 8),
    to_signed(17, 8),
    to_signed(20, 8),
    to_signed(22, 8),
    to_signed(23, 8),
    to_signed(23, 8),
    to_signed(21, 8),
    to_signed(17, 8),
    to_signed(15, 8),
    to_signed(15, 8),
    to_signed(17, 8),
    to_signed(21, 8),
    to_signed(23, 8),
    to_signed(21, 8),
    to_signed(12, 8),
    to_signed(-1, 8),
    to_signed(-11, 8),
    to_signed(-14, 8),
    to_signed(-11, 8),
    to_signed(-4, 8),
    to_signed(0, 8),
    to_signed(1, 8),
    to_signed(-2, 8),
    to_signed(-7, 8),
    to_signed(-15, 8),
    to_signed(-26, 8),
    to_signed(-33, 8),
    to_signed(-31, 8),
    to_signed(-22, 8),
    to_signed(-13, 8),
    to_signed(-8, 8),
    to_signed(-7, 8),
    to_signed(-8, 8),
    to_signed(-10, 8),
    to_signed(-12, 8),
    to_signed(-12, 8),
    to_signed(-8, 8),
    to_signed(-1, 8),
    to_signed(4, 8),
    to_signed(4, 8),
    to_signed(-2, 8),
    to_signed(-10, 8),
    to_signed(-14, 8),
    to_signed(-15, 8),
    to_signed(-11, 8),
    to_signed(-4, 8),
    to_signed(1, 8),
    to_signed(2, 8),
    to_signed(2, 8),
    to_signed(0, 8),
    to_signed(-2, 8),
    to_signed(-6, 8),
    to_signed(-10, 8),
    to_signed(-14, 8),
    to_signed(-15, 8),
    to_signed(-15, 8),
    to_signed(-14, 8),
    to_signed(-15, 8),
    to_signed(-15, 8),
    to_signed(-11, 8),
    to_signed(-3, 8),
    to_signed(4, 8),
    to_signed(7, 8),
    to_signed(7, 8),
    to_signed(9, 8),
    to_signed(13, 8),
    to_signed(15, 8),
    to_signed(14, 8),
    to_signed(13, 8),
    to_signed(12, 8),
    to_signed(10, 8),
    to_signed(10, 8),
    to_signed(10, 8),
    to_signed(10, 8),
    to_signed(9, 8),
    to_signed(9, 8),
    to_signed(9, 8),
    to_signed(8, 8),
    to_signed(6, 8),
    to_signed(4, 8),
    to_signed(-2, 8),
    to_signed(-10, 8),
    to_signed(-16, 8),
    to_signed(-19, 8),
    to_signed(-19, 8),
    to_signed(-17, 8),
    to_signed(-11, 8),
    to_signed(-2, 8),
    to_signed(7, 8),
    to_signed(11, 8),
    to_signed(15, 8),
    to_signed(20, 8),
    to_signed(22, 8),
    to_signed(19, 8),
    to_signed(16, 8),
    to_signed(15, 8),
    to_signed(17, 8),
    to_signed(21, 8),
    to_signed(27, 8),
    to_signed(32, 8),
    to_signed(33, 8),
    to_signed(31, 8),
    to_signed(30, 8),
    to_signed(29, 8),
    to_signed(26, 8),
    to_signed(21, 8),
    to_signed(14, 8),
    to_signed(1, 8),
    to_signed(-17, 8),
    to_signed(-32, 8),
    to_signed(-38, 8),
    to_signed(-36, 8),
    to_signed(-31, 8),
    to_signed(-24, 8),
    to_signed(-15, 8),
    to_signed(-10, 8),
    to_signed(-11, 8),
    to_signed(-20, 8),
    to_signed(-33, 8),
    to_signed(-45, 8),
    to_signed(-49, 8),
    to_signed(-44, 8),
    to_signed(-34, 8),
    to_signed(-23, 8),
    to_signed(-15, 8),
    to_signed(-6, 8),
    to_signed(0, 8),
    to_signed(1, 8),
    to_signed(-1, 8),
    to_signed(-1, 8),
    to_signed(1, 8),
    to_signed(0, 8),
    to_signed(-3, 8),
    to_signed(-8, 8),
    to_signed(-13, 8),
    to_signed(-16, 8),
    to_signed(-14, 8),
    to_signed(-6, 8),
    to_signed(4, 8),
    to_signed(10, 8),
    to_signed(12, 8),
    to_signed(9, 8),
    to_signed(2, 8),
    to_signed(-7, 8),
    to_signed(-12, 8),
    to_signed(-12, 8),
    to_signed(-7, 8),
    to_signed(0, 8),
    to_signed(9, 8),
    to_signed(16, 8),
    to_signed(19, 8),
    to_signed(18, 8),
    to_signed(18, 8),
    to_signed(19, 8),
    to_signed(20, 8),
    to_signed(21, 8),
    to_signed(23, 8),
    to_signed(23, 8),
    to_signed(20, 8),
    to_signed(14, 8),
    to_signed(9, 8),
    to_signed(6, 8),
    to_signed(4, 8),
    to_signed(3, 8),
    to_signed(1, 8),
    to_signed(-1, 8),
    to_signed(-4, 8),
    to_signed(-9, 8),
    to_signed(-13, 8),
    to_signed(-16, 8),
    to_signed(-18, 8),
    to_signed(-19, 8),
    to_signed(-18, 8),
    to_signed(-17, 8),
    to_signed(-18, 8),
    to_signed(-20, 8),
    to_signed(-21, 8),
    to_signed(-22, 8),
    to_signed(-20, 8),
    to_signed(-12, 8),
    to_signed(2, 8),
    to_signed(13, 8),
    to_signed(18, 8),
    to_signed(15, 8),
    to_signed(10, 8),
    to_signed(6, 8),
    to_signed(7, 8),
    to_signed(11, 8),
    to_signed(16, 8),
    to_signed(20, 8),
    to_signed(21, 8),
    to_signed(21, 8),
    to_signed(20, 8),
    to_signed(19, 8),
    to_signed(19, 8),
    to_signed(21, 8),
    to_signed(25, 8),
    to_signed(29, 8),
    to_signed(32, 8),
    to_signed(30, 8),
    to_signed(18, 8),
    to_signed(-1, 8),
    to_signed(-19, 8),
    to_signed(-26, 8),
    to_signed(-23, 8),
    to_signed(-13, 8),
    to_signed(-3, 8),
    to_signed(3, 8),
    to_signed(4, 8),
    to_signed(-2, 8),
    to_signed(-12, 8),
    to_signed(-22, 8),
    to_signed(-28, 8),
    to_signed(-30, 8),
    to_signed(-27, 8),
    to_signed(-25, 8),
    to_signed(-23, 8),
    to_signed(-23, 8),
    to_signed(-23, 8),
    to_signed(-22, 8),
    to_signed(-19, 8),
    to_signed(-15, 8),
    to_signed(-9, 8),
    to_signed(-1, 8),
    to_signed(4, 8),
    to_signed(5, 8),
    to_signed(-2, 8),
    to_signed(-14, 8),
    to_signed(-25, 8),
    to_signed(-28, 8),
    to_signed(-24, 8),
    to_signed(-16, 8),
    to_signed(-8, 8),
    to_signed(-2, 8),
    to_signed(2, 8),
    to_signed(5, 8),
    to_signed(6, 8),
    to_signed(5, 8),
    to_signed(4, 8),
    to_signed(6, 8),
    to_signed(9, 8),
    to_signed(11, 8),
    to_signed(9, 8),
    to_signed(5, 8),
    to_signed(5, 8),
    to_signed(9, 8),
    to_signed(15, 8),
    to_signed(20, 8),
    to_signed(24, 8),
    to_signed(25, 8),
    to_signed(21, 8),
    to_signed(13, 8),
    to_signed(1, 8),
    to_signed(-9, 8),
    to_signed(-12, 8),
    to_signed(-8, 8),
    to_signed(1, 8),
    to_signed(9, 8),
    to_signed(12, 8),
    to_signed(7, 8),
    to_signed(-2, 8),
    to_signed(-12, 8),
    to_signed(-18, 8),
    to_signed(-18, 8),
    to_signed(-11, 8),
    to_signed(-1, 8),
    to_signed(7, 8),
    to_signed(12, 8),
    to_signed(11, 8),
    to_signed(5, 8),
    to_signed(-3, 8),
    to_signed(-9, 8),
    to_signed(-10, 8),
    to_signed(-8, 8),
    to_signed(-3, 8),
    to_signed(1, 8),
    to_signed(4, 8),
    to_signed(4, 8),
    to_signed(3, 8),
    to_signed(0, 8),
    to_signed(-2, 8),
    to_signed(-3, 8),
    to_signed(-1, 8),
    to_signed(4, 8),
    to_signed(9, 8),
    to_signed(14, 8),
    to_signed(15, 8),
    to_signed(13, 8),
    to_signed(12, 8),
    to_signed(12, 8),
    to_signed(15, 8),
    to_signed(20, 8),
    to_signed(27, 8),
    to_signed(32, 8),
    to_signed(31, 8),
    to_signed(23, 8),
    to_signed(10, 8),
    to_signed(-8, 8),
    to_signed(-23, 8),
    to_signed(-30, 8),
    to_signed(-27, 8),
    to_signed(-19, 8),
    to_signed(-9, 8),
    to_signed(-1, 8),
    to_signed(2, 8),
    to_signed(-3, 8),
    to_signed(-14, 8),
    to_signed(-27, 8),
    to_signed(-36, 8),
    to_signed(-37, 8),
    to_signed(-31, 8),
    to_signed(-24, 8),
    to_signed(-19, 8),
    to_signed(-18, 8),
    to_signed(-19, 8),
    to_signed(-19, 8),
    to_signed(-14, 8),
    to_signed(-6, 8),
    to_signed(4, 8),
    to_signed(13, 8),
    to_signed(19, 8),
    to_signed(17, 8),
    to_signed(10, 8),
    to_signed(-1, 8),
    to_signed(-10, 8),
    to_signed(-14, 8),
    to_signed(-12, 8),
    to_signed(-6, 8),
    to_signed(1, 8),
    to_signed(6, 8),
    to_signed(9, 8),
    to_signed(12, 8),
    to_signed(14, 8),
    to_signed(17, 8),
    to_signed(16, 8),
    to_signed(13, 8),
    to_signed(8, 8),
    to_signed(2, 8),
    to_signed(-3, 8),
    to_signed(-6, 8),
    to_signed(-5, 8),
    to_signed(0, 8),
    to_signed(8, 8),
    to_signed(18, 8),
    to_signed(24, 8),
    to_signed(24, 8),
    to_signed(20, 8),
    to_signed(15, 8),
    to_signed(11, 8),
    to_signed(9, 8),
    to_signed(8, 8),
    to_signed(12, 8),
    to_signed(15, 8),
    to_signed(16, 8),
    to_signed(14, 8),
    to_signed(10, 8),
    to_signed(5, 8),
    to_signed(2, 8),
    to_signed(2, 8),
    to_signed(5, 8),
    to_signed(8, 8),
    to_signed(7, 8),
    to_signed(3, 8),
    to_signed(-3, 8),
    to_signed(-10, 8),
    to_signed(-15, 8),
    to_signed(-15, 8),
    to_signed(-13, 8),
    to_signed(-10, 8),
    to_signed(-6, 8),
    to_signed(-1, 8),
    to_signed(1, 8),
    to_signed(2, 8),
    to_signed(1, 8),
    to_signed(2, 8),
    to_signed(3, 8),
    to_signed(5, 8),
    to_signed(7, 8),
    to_signed(10, 8),
    to_signed(11, 8),
    to_signed(9, 8),
    to_signed(4, 8),
    to_signed(0, 8),
    to_signed(-2, 8),
    to_signed(0, 8),
    to_signed(7, 8),
    to_signed(15, 8),
    to_signed(21, 8),
    to_signed(23, 8),
    to_signed(21, 8),
    to_signed(15, 8),
    to_signed(7, 8),
    to_signed(0, 8),
    to_signed(-7, 8),
    to_signed(-14, 8),
    to_signed(-21, 8),
    to_signed(-22, 8),
    to_signed(-15, 8),
    to_signed(-2, 8),
    to_signed(10, 8),
    to_signed(17, 8),
    to_signed(19, 8),
    to_signed(16, 8),
    to_signed(7, 8),
    to_signed(-6, 8),
    to_signed(-20, 8),
    to_signed(-29, 8),
    to_signed(-29, 8),
    to_signed(-21, 8),
    to_signed(-9, 8),
    to_signed(2, 8),
    to_signed(7, 8),
    to_signed(9, 8),
    to_signed(9, 8),
    to_signed(7, 8),
    to_signed(6, 8),
    to_signed(9, 8),
    to_signed(13, 8),
    to_signed(14, 8),
    to_signed(12, 8),
    to_signed(7, 8),
    to_signed(0, 8),
    to_signed(-6, 8),
    to_signed(-9, 8),
    to_signed(-8, 8),
    to_signed(-4, 8),
    to_signed(0, 8),
    to_signed(1, 8),
    to_signed(-2, 8),
    to_signed(-8, 8),
    to_signed(-14, 8),
    to_signed(-17, 8),
    to_signed(-18, 8),
    to_signed(-19, 8),
    to_signed(-19, 8),
    to_signed(-19, 8),
    to_signed(-19, 8),
    to_signed(-19, 8),
    to_signed(-16, 8),
    to_signed(-10, 8),
    to_signed(-3, 8),
    to_signed(4, 8),
    to_signed(9, 8),
    to_signed(11, 8),
    to_signed(8, 8),
    to_signed(3, 8),
    to_signed(2, 8),
    to_signed(4, 8),
    to_signed(9, 8),
    to_signed(12, 8),
    to_signed(12, 8),
    to_signed(8, 8),
    to_signed(1, 8),
    to_signed(-6, 8),
    to_signed(-10, 8),
    to_signed(-10, 8),
    to_signed(-6, 8),
    to_signed(0, 8),
    to_signed(5, 8),
    to_signed(6, 8),
    to_signed(0, 8),
    to_signed(-8, 8),
    to_signed(-14, 8),
    to_signed(-15, 8),
    to_signed(-13, 8),
    to_signed(-8, 8),
    to_signed(-3, 8),
    to_signed(2, 8),
    to_signed(5, 8),
    to_signed(5, 8),
    to_signed(4, 8),
    to_signed(2, 8),
    to_signed(2, 8),
    to_signed(3, 8),
    to_signed(3, 8),
    to_signed(1, 8),
    to_signed(0, 8),
    to_signed(0, 8),
    to_signed(0, 8),
    to_signed(-1, 8),
    to_signed(-3, 8),
    to_signed(-1, 8),
    to_signed(4, 8),
    to_signed(9, 8),
    to_signed(12, 8),
    to_signed(13, 8),
    to_signed(14, 8),
    to_signed(14, 8),
    to_signed(15, 8),
    to_signed(17, 8),
    to_signed(20, 8),
    to_signed(18, 8),
    to_signed(10, 8),
    to_signed(-2, 8),
    to_signed(-16, 8),
    to_signed(-24, 8),
    to_signed(-24, 8),
    to_signed(-15, 8),
    to_signed(-4, 8),
    to_signed(2, 8),
    to_signed(3, 8),
    to_signed(0, 8),
    to_signed(-8, 8),
    to_signed(-22, 8),
    to_signed(-36, 8),
    to_signed(-44, 8),
    to_signed(-44, 8),
    to_signed(-38, 8),
    to_signed(-28, 8),
    to_signed(-18, 8),
    to_signed(-14, 8),
    to_signed(-15, 8),
    to_signed(-17, 8),
    to_signed(-15, 8),
    to_signed(-10, 8),
    to_signed(-3, 8),
    to_signed(2, 8),
    to_signed(3, 8),
    to_signed(-2, 8),
    to_signed(-12, 8),
    to_signed(-21, 8),
    to_signed(-25, 8),
    to_signed(-22, 8),
    to_signed(-13, 8),
    to_signed(-2, 8),
    to_signed(6, 8),
    to_signed(8, 8),
    to_signed(7, 8),
    to_signed(4, 8),
    to_signed(1, 8),
    to_signed(-2, 8),
    to_signed(-4, 8),
    to_signed(-3, 8),
    to_signed(-3, 8),
    to_signed(-2, 8),
    to_signed(-1, 8),
    to_signed(2, 8),
    to_signed(4, 8),
    to_signed(6, 8),
    to_signed(6, 8),
    to_signed(6, 8),
    to_signed(5, 8),
    to_signed(3, 8),
    to_signed(1, 8),
    to_signed(0, 8),
    to_signed(0, 8),
    to_signed(1, 8),
    to_signed(1, 8),
    to_signed(-1, 8),
    to_signed(-5, 8),
    to_signed(-10, 8),
    to_signed(-13, 8),
    to_signed(-14, 8),
    to_signed(-13, 8),
    to_signed(-11, 8),
    to_signed(-7, 8),
    to_signed(-3, 8),
    to_signed(-4, 8),
    to_signed(-10, 8),
    to_signed(-18, 8),
    to_signed(-24, 8),
    to_signed(-28, 8),
    to_signed(-29, 8),
    to_signed(-28, 8),
    to_signed(-25, 8),
    to_signed(-19, 8),
    to_signed(-13, 8),
    to_signed(-9, 8),
    to_signed(-8, 8),
    to_signed(-7, 8),
    to_signed(-7, 8),
    to_signed(-4, 8),
    to_signed(2, 8),
    to_signed(7, 8),
    to_signed(8, 8),
    to_signed(6, 8),
    to_signed(5, 8),
    to_signed(5, 8),
    to_signed(8, 8),
    to_signed(14, 8),
    to_signed(22, 8),
    to_signed(29, 8),
    to_signed(35, 8),
    to_signed(37, 8),
    to_signed(37, 8),
    to_signed(34, 8),
    to_signed(28, 8),
    to_signed(20, 8),
    to_signed(14, 8),
    to_signed(14, 8),
    to_signed(20, 8),
    to_signed(29, 8),
    to_signed(33, 8),
    to_signed(28, 8),
    to_signed(14, 8),
    to_signed(-2, 8),
    to_signed(-14, 8),
    to_signed(-16, 8),
    to_signed(-12, 8),
    to_signed(-3, 8),
    to_signed(2, 8),
    to_signed(1, 8),
    to_signed(-7, 8),
    to_signed(-20, 8),
    to_signed(-32, 8),
    to_signed(-41, 8),
    to_signed(-44, 8),
    to_signed(-40, 8),
    to_signed(-32, 8),
    to_signed(-24, 8),
    to_signed(-20, 8),
    to_signed(-20, 8),
    to_signed(-24, 8),
    to_signed(-27, 8),
    to_signed(-26, 8),
    to_signed(-16, 8),
    to_signed(-4, 8),
    to_signed(5, 8),
    to_signed(8, 8),
    to_signed(4, 8),
    to_signed(-4, 8),
    to_signed(-12, 8),
    to_signed(-13, 8),
    to_signed(-6, 8),
    to_signed(4, 8),
    to_signed(13, 8),
    to_signed(15, 8),
    to_signed(13, 8),
    to_signed(7, 8),
    to_signed(2, 8),
    to_signed(-2, 8),
    to_signed(-2, 8),
    to_signed(-1, 8),
    to_signed(1, 8),
    to_signed(3, 8),
    to_signed(4, 8),
    to_signed(4, 8),
    to_signed(5, 8),
    to_signed(7, 8),
    to_signed(11, 8),
    to_signed(14, 8),
    to_signed(13, 8),
    to_signed(9, 8),
    to_signed(4, 8),
    to_signed(2, 8),
    to_signed(3, 8),
    to_signed(6, 8),
    to_signed(9, 8),
    to_signed(10, 8),
    to_signed(9, 8),
    to_signed(7, 8),
    to_signed(3, 8),
    to_signed(-2, 8),
    to_signed(-7, 8),
    to_signed(-10, 8),
    to_signed(-12, 8),
    to_signed(-13, 8),
    to_signed(-15, 8),
    to_signed(-16, 8),
    to_signed(-16, 8),
    to_signed(-14, 8),
    to_signed(-11, 8),
    to_signed(-8, 8),
    to_signed(-7, 8),
    to_signed(-9, 8),
    to_signed(-14, 8),
    to_signed(-16, 8),
    to_signed(-17, 8),
    to_signed(-15, 8),
    to_signed(-13, 8),
    to_signed(-10, 8),
    to_signed(-8, 8),
    to_signed(-7, 8),
    to_signed(-6, 8),
    to_signed(-4, 8),
    to_signed(-2, 8),
    to_signed(0, 8),
    to_signed(1, 8),
    to_signed(1, 8),
    to_signed(0, 8),
    to_signed(-1, 8),
    to_signed(0, 8),
    to_signed(4, 8),
    to_signed(10, 8),
    to_signed(16, 8),
    to_signed(21, 8),
    to_signed(22, 8),
    to_signed(20, 8),
    to_signed(16, 8),
    to_signed(13, 8),
    to_signed(12, 8),
    to_signed(14, 8),
    to_signed(18, 8),
    to_signed(23, 8),
    to_signed(26, 8),
    to_signed(21, 8),
    to_signed(10, 8),
    to_signed(-2, 8),
    to_signed(-10, 8),
    to_signed(-11, 8),
    to_signed(-7, 8),
    to_signed(-2, 8),
    to_signed(0, 8),
    to_signed(-1, 8),
    to_signed(-5, 8),
    to_signed(-11, 8),
    to_signed(-19, 8),
    to_signed(-26, 8),
    to_signed(-27, 8),
    to_signed(-24, 8),
    to_signed(-20, 8),
    to_signed(-19, 8),
    to_signed(-20, 8),
    to_signed(-22, 8),
    to_signed(-23, 8),
    to_signed(-21, 8),
    to_signed(-16, 8),
    to_signed(-10, 8),
    to_signed(-4, 8),
    to_signed(1, 8),
    to_signed(1, 8),
    to_signed(-3, 8),
    to_signed(-8, 8),
    to_signed(-11, 8),
    to_signed(-10, 8),
    to_signed(-4, 8),
    to_signed(4, 8),
    to_signed(12, 8),
    to_signed(16, 8),
    to_signed(15, 8),
    to_signed(12, 8),
    to_signed(9, 8),
    to_signed(7, 8),
    to_signed(8, 8),
    to_signed(10, 8),
    to_signed(13, 8),
    to_signed(14, 8),
    to_signed(12, 8),
    to_signed(8, 8),
    to_signed(4, 8),
    to_signed(3, 8),
    to_signed(8, 8),
    to_signed(16, 8),
    to_signed(22, 8),
    to_signed(22, 8),
    to_signed(20, 8),
    to_signed(16, 8),
    to_signed(13, 8),
    to_signed(12, 8),
    to_signed(14, 8),
    to_signed(16, 8),
    to_signed(17, 8),
    to_signed(17, 8),
    to_signed(14, 8),
    to_signed(10, 8),
    to_signed(3, 8),
    to_signed(-4, 8),
    to_signed(-9, 8),
    to_signed(-12, 8),
    to_signed(-11, 8),
    to_signed(-8, 8),
    to_signed(-6, 8),
    to_signed(-6, 8),
    to_signed(-10, 8),
    to_signed(-13, 8),
    to_signed(-16, 8),
    to_signed(-18, 8),
    to_signed(-19, 8),
    to_signed(-16, 8),
    to_signed(-10, 8),
    to_signed(-4, 8),
    to_signed(0, 8),
    to_signed(2, 8),
    to_signed(2, 8),
    to_signed(2, 8),
    to_signed(3, 8),
    to_signed(3, 8),
    to_signed(4, 8),
    to_signed(3, 8),
    to_signed(2, 8),
    to_signed(0, 8),
    to_signed(-2, 8),
    to_signed(-3, 8),
    to_signed(-2, 8),
    to_signed(0, 8),
    to_signed(3, 8),
    to_signed(6, 8),
    to_signed(8, 8),
    to_signed(10, 8),
    to_signed(9, 8),
    to_signed(6, 8),
    to_signed(4, 8),
    to_signed(6, 8),
    to_signed(11, 8),
    to_signed(17, 8),
    to_signed(22, 8),
    to_signed(26, 8),
    to_signed(29, 8),
    to_signed(28, 8),
    to_signed(22, 8),
    to_signed(15, 8),
    to_signed(7, 8),
    to_signed(3, 8),
    to_signed(1, 8),
    to_signed(1, 8),
    to_signed(2, 8),
    to_signed(4, 8),
    to_signed(3, 8),
    to_signed(-1, 8),
    to_signed(-7, 8),
    to_signed(-14, 8),
    to_signed(-19, 8),
    to_signed(-21, 8),
    to_signed(-22, 8),
    to_signed(-21, 8),
    to_signed(-21, 8),
    to_signed(-19, 8),
    to_signed(-18, 8),
    to_signed(-18, 8),
    to_signed(-19, 8),
    to_signed(-16, 8),
    to_signed(-11, 8),
    to_signed(-6, 8),
    to_signed(-2, 8),
    to_signed(-1, 8),
    to_signed(-5, 8),
    to_signed(-10, 8),
    to_signed(-13, 8),
    to_signed(-12, 8),
    to_signed(-5, 8),
    to_signed(1, 8),
    to_signed(4, 8),
    to_signed(4, 8),
    to_signed(3, 8),
    to_signed(1, 8),
    to_signed(1, 8),
    to_signed(2, 8),
    to_signed(5, 8),
    to_signed(7, 8),
    to_signed(9, 8),
    to_signed(10, 8),
    to_signed(9, 8),
    to_signed(6, 8),
    to_signed(5, 8),
    to_signed(7, 8),
    to_signed(10, 8),
    to_signed(11, 8),
    to_signed(11, 8),
    to_signed(10, 8),
    to_signed(8, 8),
    to_signed(4, 8),
    to_signed(1, 8),
    to_signed(2, 8),
    to_signed(6, 8),
    to_signed(9, 8),
    to_signed(11, 8),
    to_signed(10, 8),
    to_signed(6, 8),
    to_signed(0, 8),
    to_signed(-6, 8),
    to_signed(-11, 8),
    to_signed(-12, 8),
    to_signed(-9, 8),
    to_signed(-2, 8),
    to_signed(3, 8),
    to_signed(4, 8),
    to_signed(0, 8),
    to_signed(-6, 8),
    to_signed(-14, 8),
    to_signed(-21, 8),
    to_signed(-26, 8),
    to_signed(-25, 8),
    to_signed(-21, 8),
    to_signed(-15, 8),
    to_signed(-11, 8),
    to_signed(-9, 8),
    to_signed(-9, 8),
    to_signed(-11, 8),
    to_signed(-13, 8),
    to_signed(-12, 8),
    to_signed(-11, 8),
    to_signed(-11, 8),
    to_signed(-11, 8),
    to_signed(-11, 8),
    to_signed(-10, 8),
    to_signed(-9, 8),
    to_signed(-7, 8),
    to_signed(-3, 8),
    to_signed(2, 8),
    to_signed(8, 8),
    to_signed(12, 8),
    to_signed(13, 8),
    to_signed(12, 8),
    to_signed(9, 8),
    to_signed(7, 8),
    to_signed(8, 8),
    to_signed(11, 8),
    to_signed(12, 8),
    to_signed(13, 8),
    to_signed(17, 8),
    to_signed(22, 8),
    to_signed(26, 8),
    to_signed(27, 8),
    to_signed(28, 8),
    to_signed(28, 8),
    to_signed(25, 8),
    to_signed(18, 8),
    to_signed(9, 8),
    to_signed(2, 8),
    to_signed(-1, 8),
    to_signed(-1, 8),
    to_signed(0, 8),
    to_signed(-2, 8),
    to_signed(-4, 8),
    to_signed(-6, 8),
    to_signed(-9, 8),
    to_signed(-13, 8),
    to_signed(-19, 8),
    to_signed(-24, 8),
    to_signed(-26, 8),
    to_signed(-27, 8),
    to_signed(-27, 8),
    to_signed(-29, 8),
    to_signed(-31, 8),
    to_signed(-32, 8),
    to_signed(-30, 8),
    to_signed(-25, 8),
    to_signed(-19, 8),
    to_signed(-15, 8),
    to_signed(-13, 8),
    to_signed(-13, 8),
    to_signed(-13, 8),
    to_signed(-14, 8),
    to_signed(-16, 8),
    to_signed(-18, 8),
    to_signed(-17, 8),
    to_signed(-13, 8),
    to_signed(-8, 8),
    to_signed(-2, 8),
    to_signed(1, 8),
    to_signed(2, 8),
    to_signed(2, 8),
    to_signed(2, 8),
    to_signed(4, 8),
    to_signed(5, 8),
    to_signed(6, 8),
    to_signed(8, 8),
    to_signed(10, 8),
    to_signed(12, 8),
    to_signed(12, 8),
    to_signed(12, 8),
    to_signed(14, 8),
    to_signed(17, 8),
    to_signed(20, 8),
    to_signed(23, 8),
    to_signed(25, 8),
    to_signed(24, 8),
    to_signed(20, 8),
    to_signed(17, 8),
    to_signed(14, 8),
    to_signed(13, 8),
    to_signed(13, 8),
    to_signed(12, 8),
    to_signed(11, 8),
    to_signed(9, 8),
    to_signed(6, 8),
    to_signed(2, 8),
    to_signed(-2, 8),
    to_signed(-6, 8),
    to_signed(-8, 8),
    to_signed(-9, 8),
    to_signed(-9, 8),
    to_signed(-10, 8),
    to_signed(-11, 8),
    to_signed(-13, 8),
    to_signed(-17, 8),
    to_signed(-22, 8),
    to_signed(-26, 8),
    to_signed(-28, 8),
    to_signed(-28, 8),
    to_signed(-26, 8),
    to_signed(-22, 8),
    to_signed(-18, 8),
    to_signed(-15, 8),
    to_signed(-14, 8),
    to_signed(-15, 8),
    to_signed(-14, 8),
    to_signed(-13, 8),
    to_signed(-14, 8),
    to_signed(-15, 8),
    to_signed(-12, 8),
    to_signed(-9, 8),
    to_signed(-6, 8),
    to_signed(-5, 8),
    to_signed(-2, 8),
    to_signed(3, 8),
    to_signed(9, 8),
    to_signed(14, 8),
    to_signed(16, 8),
    to_signed(15, 8),
    to_signed(12, 8),
    to_signed(11, 8),
    to_signed(13, 8),
    to_signed(15, 8),
    to_signed(17, 8),
    to_signed(21, 8),
    to_signed(26, 8),
    to_signed(29, 8),
    to_signed(28, 8),
    to_signed(26, 8),
    to_signed(24, 8),
    to_signed(23, 8),
    to_signed(24, 8),
    to_signed(25, 8),
    to_signed(25, 8),
    to_signed(22, 8),
    to_signed(18, 8),
    to_signed(13, 8),
    to_signed(10, 8),
    to_signed(8, 8),
    to_signed(7, 8),
    to_signed(6, 8),
    to_signed(4, 8),
    to_signed(1, 8),
    to_signed(-3, 8),
    to_signed(-9, 8),
    to_signed(-13, 8),
    to_signed(-16, 8),
    to_signed(-17, 8),
    to_signed(-17, 8),
    to_signed(-16, 8),
    to_signed(-17, 8),
    to_signed(-20, 8),
    to_signed(-23, 8),
    to_signed(-25, 8),
    to_signed(-25, 8),
    to_signed(-23, 8),
    to_signed(-19, 8),
    to_signed(-15, 8),
    to_signed(-13, 8),
    to_signed(-12, 8),
    to_signed(-10, 8),
    to_signed(-8, 8),
    to_signed(-8, 8),
    to_signed(-12, 8),
    to_signed(-14, 8),
    to_signed(-13, 8),
    to_signed(-9, 8),
    to_signed(-4, 8),
    to_signed(-1, 8),
    to_signed(0, 8),
    to_signed(-1, 8),
    to_signed(-2, 8),
    to_signed(-3, 8),
    to_signed(-3, 8),
    to_signed(-3, 8),
    to_signed(-2, 8),
    to_signed(0, 8),
    to_signed(2, 8),
    to_signed(5, 8),
    to_signed(9, 8),
    to_signed(12, 8),
    to_signed(14, 8),
    to_signed(16, 8),
    to_signed(18, 8),
    to_signed(21, 8),
    to_signed(23, 8),
    to_signed(24, 8),
    to_signed(23, 8),
    to_signed(21, 8),
    to_signed(20, 8),
    to_signed(20, 8),
    to_signed(19, 8),
    to_signed(17, 8),
    to_signed(15, 8),
    to_signed(14, 8),
    to_signed(13, 8),
    to_signed(13, 8),
    to_signed(13, 8),
    to_signed(11, 8),
    to_signed(6, 8),
    to_signed(1, 8),
    to_signed(-1, 8),
    to_signed(-3, 8),
    to_signed(-4, 8),
    to_signed(-4, 8),
    to_signed(-3, 8),
    to_signed(-4, 8),
    to_signed(-6, 8),
    to_signed(-6, 8),
    to_signed(-8, 8),
    to_signed(-11, 8),
    to_signed(-13, 8),
    to_signed(-12, 8),
    to_signed(-10, 8),
    to_signed(-7, 8),
    to_signed(-5, 8),
    to_signed(-4, 8),
    to_signed(-6, 8),
    to_signed(-8, 8),
    to_signed(-9, 8),
    to_signed(-9, 8),
    to_signed(-8, 8),
    to_signed(-6, 8),
    to_signed(-3, 8),
    to_signed(-1, 8),
    to_signed(-1, 8),
    to_signed(-2, 8),
    to_signed(-1, 8),
    to_signed(1, 8),
    to_signed(3, 8),
    to_signed(5, 8),
    to_signed(8, 8),
    to_signed(9, 8),
    to_signed(9, 8),
    to_signed(10, 8),
    to_signed(11, 8),
    to_signed(13, 8),
    to_signed(14, 8),
    to_signed(15, 8),
    to_signed(17, 8),
    to_signed(20, 8),
    to_signed(23, 8),
    to_signed(24, 8),
    to_signed(24, 8),
    to_signed(24, 8),
    to_signed(24, 8),
    to_signed(22, 8),
    to_signed(20, 8),
    to_signed(18, 8),
    to_signed(19, 8),
    to_signed(19, 8),
    to_signed(18, 8),
    to_signed(17, 8),
    to_signed(17, 8),
    to_signed(15, 8),
    to_signed(11, 8),
    to_signed(7, 8),
    to_signed(4, 8),
    to_signed(1, 8),
    to_signed(1, 8),
    to_signed(0, 8),
    to_signed(-3, 8),
    to_signed(-8, 8),
    to_signed(-11, 8),
    to_signed(-13, 8),
    to_signed(-15, 8),
    to_signed(-16, 8),
    to_signed(-17, 8),
    to_signed(-15, 8),
    to_signed(-14, 8),
    to_signed(-14, 8),
    to_signed(-17, 8),
    to_signed(-20, 8),
    to_signed(-21, 8),
    to_signed(-20, 8),
    to_signed(-16, 8),
    to_signed(-11, 8),
    to_signed(-9, 8),
    to_signed(-7, 8),
    to_signed(-8, 8),
    to_signed(-10, 8),
    to_signed(-11, 8),
    to_signed(-10, 8),
    to_signed(-5, 8),
    to_signed(-2, 8),
    to_signed(1, 8),
    to_signed(1, 8),
    to_signed(2, 8),
    to_signed(1, 8),
    to_signed(2, 8),
    to_signed(4, 8),
    to_signed(7, 8),
    to_signed(10, 8),
    to_signed(12, 8),
    to_signed(13, 8),
    to_signed(14, 8),
    to_signed(14, 8),
    to_signed(14, 8),
    to_signed(13, 8),
    to_signed(12, 8),
    to_signed(13, 8),
    to_signed(13, 8),
    to_signed(12, 8),
    to_signed(9, 8),
    to_signed(8, 8),
    to_signed(6, 8),
    to_signed(6, 8),
    to_signed(6, 8),
    to_signed(7, 8),
    to_signed(6, 8),
    to_signed(2, 8),
    to_signed(-1, 8),
    to_signed(-4, 8),
    to_signed(-8, 8),
    to_signed(-12, 8),
    to_signed(-12, 8),
    to_signed(-11, 8),
    to_signed(-10, 8),
    to_signed(-9, 8),
    to_signed(-8, 8),
    to_signed(-9, 8),
    to_signed(-10, 8),
    to_signed(-12, 8),
    to_signed(-15, 8),
    to_signed(-18, 8),
    to_signed(-20, 8),
    to_signed(-19, 8),
    to_signed(-17, 8),
    to_signed(-15, 8),
    to_signed(-12, 8),
    to_signed(-10, 8),
    to_signed(-9, 8),
    to_signed(-11, 8),
    to_signed(-13, 8),
    to_signed(-15, 8),
    to_signed(-14, 8),
    to_signed(-12, 8),
    to_signed(-8, 8),
    to_signed(-5, 8),
    to_signed(-4, 8),
    to_signed(-4, 8),
    to_signed(-4, 8),
    to_signed(-3, 8),
    to_signed(-1, 8),
    to_signed(0, 8),
    to_signed(1, 8),
    to_signed(1, 8),
    to_signed(1, 8),
    to_signed(2, 8),
    to_signed(3, 8),
    to_signed(5, 8),
    to_signed(7, 8),
    to_signed(10, 8),
    to_signed(13, 8),
    to_signed(15, 8),
    to_signed(15, 8),
    to_signed(13, 8),
    to_signed(12, 8),
    to_signed(12, 8),
    to_signed(13, 8),
    to_signed(13, 8),
    to_signed(13, 8),
    to_signed(12, 8),
    to_signed(12, 8),
    to_signed(11, 8),
    to_signed(7, 8),
    to_signed(3, 8),
    to_signed(0, 8),
    to_signed(-2, 8),
    to_signed(-4, 8),
    to_signed(-6, 8),
    to_signed(-8, 8),
    to_signed(-11, 8),
    to_signed(-14, 8),
    to_signed(-17, 8),
    to_signed(-18, 8),
    to_signed(-18, 8),
    to_signed(-16, 8),
    to_signed(-14, 8),
    to_signed(-13, 8),
    to_signed(-15, 8),
    to_signed(-17, 8),
    to_signed(-18, 8),
    to_signed(-18, 8),
    to_signed(-18, 8),
    to_signed(-15, 8),
    to_signed(-12, 8),
    to_signed(-10, 8),
    to_signed(-11, 8),
    to_signed(-12, 8),
    to_signed(-13, 8),
    to_signed(-14, 8),
    to_signed(-14, 8),
    to_signed(-14, 8),
    to_signed(-12, 8),
    to_signed(-10, 8),
    to_signed(-7, 8),
    to_signed(-4, 8),
    to_signed(-3, 8),
    to_signed(-3, 8),
    to_signed(-4, 8),
    to_signed(-4, 8),
    to_signed(-4, 8),
    to_signed(-2, 8),
    to_signed(1, 8),
    to_signed(2, 8),
    to_signed(3, 8),
    to_signed(4, 8),
    to_signed(6, 8),
    to_signed(8, 8),
    to_signed(8, 8),
    to_signed(8, 8),
    to_signed(7, 8),
    to_signed(6, 8),
    to_signed(4, 8),
    to_signed(3, 8),
    to_signed(1, 8),
    to_signed(0, 8),
    to_signed(-1, 8),
    to_signed(0, 8),
    to_signed(1, 8),
    to_signed(3, 8),
    to_signed(5, 8),
    to_signed(5, 8),
    to_signed(3, 8),
    to_signed(1, 8),
    to_signed(-1, 8),
    to_signed(-2, 8),
    to_signed(-2, 8),
    to_signed(-2, 8),
    to_signed(-3, 8),
    to_signed(-4, 8),
    to_signed(-6, 8),
    to_signed(-8, 8),
    to_signed(-9, 8),
    to_signed(-9, 8),
    to_signed(-9, 8),
    to_signed(-9, 8),
    to_signed(-10, 8),
    to_signed(-11, 8),
    to_signed(-13, 8),
    to_signed(-13, 8),
    to_signed(-12, 8),
    to_signed(-10, 8),
    to_signed(-8, 8),
    to_signed(-6, 8),
    to_signed(-5, 8),
    to_signed(-5, 8),
    to_signed(-4, 8),
    to_signed(-5, 8),
    to_signed(-7, 8),
    to_signed(-6, 8),
    to_signed(-3, 8),
    to_signed(0, 8),
    to_signed(2, 8),
    to_signed(2, 8),
    to_signed(2, 8),
    to_signed(2, 8),
    to_signed(3, 8),
    to_signed(4, 8),
    to_signed(5, 8),
    to_signed(5, 8),
    to_signed(5, 8),
    to_signed(4, 8),
    to_signed(4, 8),
    to_signed(5, 8),
    to_signed(7, 8),
    to_signed(8, 8),
    to_signed(9, 8),
    to_signed(11, 8),
    to_signed(14, 8),
    to_signed(16, 8),
    to_signed(15, 8),
    to_signed(14, 8),
    to_signed(13, 8),
    to_signed(12, 8),
    to_signed(11, 8),
    to_signed(10, 8),
    to_signed(8, 8),
    to_signed(6, 8),
    to_signed(5, 8),
    to_signed(4, 8),
    to_signed(3, 8),
    to_signed(3, 8),
    to_signed(3, 8),
    to_signed(3, 8),
    to_signed(2, 8),
    to_signed(1, 8),
    to_signed(0, 8),
    to_signed(-1, 8),
    to_signed(-3, 8),
    to_signed(-5, 8),
    to_signed(-6, 8),
    to_signed(-5, 8),
    to_signed(-4, 8),
    to_signed(-4, 8),
    to_signed(-4, 8),
    to_signed(-4, 8),
    to_signed(-5, 8),
    to_signed(-7, 8),
    to_signed(-9, 8),
    to_signed(-10, 8),
    to_signed(-10, 8),
    to_signed(-9, 8),
    to_signed(-7, 8),
    to_signed(-7, 8),
    to_signed(-7, 8),
    to_signed(-8, 8),
    to_signed(-8, 8),
    to_signed(-8, 8),
    to_signed(-7, 8),
    to_signed(-5, 8),
    to_signed(-2, 8),
    to_signed(0, 8),
    to_signed(1, 8),
    to_signed(2, 8),
    to_signed(1, 8),
    to_signed(1, 8),
    to_signed(1, 8),
    to_signed(1, 8),
    to_signed(1, 8),
    to_signed(2, 8),
    to_signed(2, 8),
    to_signed(1, 8),
    to_signed(0, 8),
    to_signed(1, 8),
    to_signed(2, 8),
    to_signed(3, 8),
    to_signed(3, 8),
    to_signed(3, 8),
    to_signed(2, 8),
    to_signed(1, 8),
    to_signed(0, 8),
    to_signed(0, 8),
    to_signed(-1, 8),
    to_signed(-2, 8),
    to_signed(-1, 8),
    to_signed(0, 8),
    to_signed(1, 8),
    to_signed(0, 8),
    to_signed(0, 8),
    to_signed(-2, 8),
    to_signed(-4, 8),
    to_signed(-7, 8),
    to_signed(-8, 8),
    to_signed(-9, 8),
    to_signed(-9, 8),
    to_signed(-9, 8),
    to_signed(-10, 8),
    to_signed(-10, 8),
    to_signed(-12, 8),
    to_signed(-12, 8),
    to_signed(-13, 8),
    to_signed(-12, 8),
    to_signed(-11, 8),
    to_signed(-9, 8),
    to_signed(-7, 8),
    to_signed(-6, 8),
    to_signed(-6, 8),
    to_signed(-6, 8),
    to_signed(-7, 8),
    to_signed(-7, 8),
    to_signed(-7, 8),
    to_signed(-7, 8),
    to_signed(-8, 8),
    to_signed(-8, 8),
    to_signed(-8, 8),
    to_signed(-7, 8),
    to_signed(-6, 8),
    to_signed(-5, 8),
    to_signed(-5, 8),
    to_signed(-5, 8),
    to_signed(-5, 8),
    to_signed(-5, 8),
    to_signed(-4, 8),
    to_signed(-2, 8),
    to_signed(1, 8),
    to_signed(2, 8),
    to_signed(3, 8),
    to_signed(4, 8),
    to_signed(6, 8),
    to_signed(7, 8),
    to_signed(7, 8),
    to_signed(7, 8),
    to_signed(7, 8),
    to_signed(7, 8),
    to_signed(6, 8),
    to_signed(4, 8),
    to_signed(1, 8),
    to_signed(-1, 8),
    to_signed(-1, 8),
    to_signed(0, 8),
    to_signed(0, 8),
    to_signed(1, 8),
    to_signed(1, 8),
    to_signed(1, 8),
    to_signed(1, 8),
    to_signed(0, 8),
    to_signed(0, 8),
    to_signed(0, 8),
    to_signed(0, 8),
    to_signed(0, 8),
    to_signed(1, 8),
    to_signed(2, 8),
    to_signed(2, 8),
    to_signed(2, 8),
    to_signed(2, 8),
    to_signed(2, 8),
    to_signed(2, 8),
    to_signed(1, 8),
    to_signed(1, 8),
    to_signed(0, 8),
    to_signed(-1, 8),
    to_signed(-1, 8),
    to_signed(-1, 8),
    to_signed(-1, 8),
    to_signed(0, 8),
    to_signed(0, 8),
    to_signed(0, 8),
    to_signed(0, 8),
    to_signed(0, 8),
    to_signed(1, 8),
    to_signed(2, 8),
    to_signed(4, 8),
    to_signed(6, 8),
    to_signed(7, 8),
    to_signed(7, 8),
    to_signed(7, 8),
    to_signed(7, 8),
    to_signed(6, 8),
    to_signed(5, 8),
    to_signed(3, 8),
    to_signed(3, 8),
    to_signed(4, 8),
    to_signed(4, 8),
    to_signed(4, 8),
    to_signed(4, 8),
    to_signed(4, 8),
    to_signed(2, 8),
    to_signed(1, 8),
    to_signed(-1, 8),
    to_signed(-1, 8),
    to_signed(0, 8),
    to_signed(2, 8),
    to_signed(3, 8),
    to_signed(3, 8),
    to_signed(4, 8),
    to_signed(4, 8),
    to_signed(4, 8),
    to_signed(4, 8),
    to_signed(3, 8),
    to_signed(2, 8),
    to_signed(1, 8),
    to_signed(0, 8),
    to_signed(-1, 8),
    to_signed(-2, 8),
    to_signed(-2, 8),
    to_signed(-2, 8),
    to_signed(-2, 8),
    to_signed(-3, 8),
    to_signed(-3, 8),
    to_signed(-4, 8),
    to_signed(-6, 8),
    to_signed(-8, 8),
    to_signed(-8, 8),
    to_signed(-9, 8),
    to_signed(-9, 8),
    to_signed(-8, 8),
    to_signed(-7, 8),
    to_signed(-6, 8),
    to_signed(-6, 8),
    to_signed(-7, 8),
    to_signed(-8, 8),
    to_signed(-8, 8),
    to_signed(-7, 8),
    to_signed(-7, 8),
    to_signed(-7, 8),
    to_signed(-7, 8),
    to_signed(-6, 8),
    to_signed(-6, 8),
    to_signed(-7, 8),
    to_signed(-8, 8),
    to_signed(-9, 8),
    to_signed(-8, 8),
    to_signed(-7, 8),
    to_signed(-6, 8),
    to_signed(-4, 8),
    to_signed(-3, 8),
    to_signed(-2, 8),
    to_signed(0, 8),
    to_signed(1, 8),
    to_signed(1, 8),
    to_signed(2, 8),
    to_signed(2, 8),
    to_signed(1, 8),
    to_signed(0, 8),
    to_signed(0, 8),
    to_signed(-1, 8),
    to_signed(-3, 8),
    to_signed(-3, 8),
    to_signed(-2, 8),
    to_signed(-1, 8),
    to_signed(-1, 8),
    to_signed(-2, 8),
    to_signed(-2, 8),
    to_signed(-3, 8),
    to_signed(-4, 8),
    to_signed(-4, 8),
    to_signed(-4, 8),
    to_signed(-3, 8),
    to_signed(-4, 8),
    to_signed(-4, 8),
    to_signed(-4, 8),
    to_signed(-4, 8),
    to_signed(-3, 8),
    to_signed(-2, 8),
    to_signed(-2, 8),
    to_signed(-2, 8),
    to_signed(-3, 8),
    to_signed(-4, 8),
    to_signed(-4, 8),
    to_signed(-3, 8),
    to_signed(-1, 8),
    to_signed(0, 8),
    to_signed(0, 8),
    to_signed(-1, 8),
    to_signed(-2, 8),
    to_signed(-3, 8),
    to_signed(-3, 8),
    to_signed(-3, 8),
    to_signed(-2, 8),
    to_signed(1, 8),
    to_signed(4, 8),
    to_signed(6, 8),
    to_signed(6, 8),
    to_signed(6, 8),
    to_signed(6, 8),
    to_signed(5, 8),
    to_signed(4, 8),
    to_signed(3, 8),
    to_signed(4, 8),
    to_signed(4, 8),
    to_signed(4, 8),
    to_signed(5, 8),
    to_signed(6, 8),
    to_signed(7, 8),
    to_signed(6, 8),
    to_signed(4, 8),
    to_signed(1, 8),
    to_signed(-1, 8),
    to_signed(-2, 8),
    to_signed(-1, 8),
    to_signed(0, 8),
    to_signed(1, 8),
    to_signed(2, 8),
    to_signed(2, 8),
    to_signed(2, 8),
    to_signed(1, 8),
    to_signed(-1, 8),
    to_signed(-2, 8),
    to_signed(-2, 8),
    to_signed(-3, 8),
    to_signed(-3, 8),
    to_signed(-3, 8),
    to_signed(-3, 8),
    to_signed(-3, 8),
    to_signed(-3, 8),
    to_signed(-4, 8),
    to_signed(-5, 8),
    to_signed(-6, 8),
    to_signed(-7, 8),
    to_signed(-8, 8),
    to_signed(-8, 8),
    to_signed(-8, 8),
    to_signed(-7, 8),
    to_signed(-6, 8),
    to_signed(-5, 8),
    to_signed(-3, 8),
    to_signed(-1, 8),
    to_signed(1, 8),
    to_signed(1, 8),
    to_signed(2, 8),
    to_signed(2, 8),
    to_signed(3, 8),
    to_signed(3, 8),
    to_signed(3, 8),
    to_signed(3, 8),
    to_signed(5, 8),
    to_signed(6, 8),
    to_signed(6, 8),
    to_signed(4, 8),
    to_signed(2, 8),
    to_signed(0, 8),
    to_signed(0, 8),
    to_signed(0, 8),
    to_signed(1, 8),
    to_signed(2, 8),
    to_signed(3, 8),
    to_signed(4, 8),
    to_signed(4, 8),
    to_signed(3, 8),
    to_signed(3, 8),
    to_signed(2, 8),
    to_signed(1, 8),
    to_signed(1, 8),
    to_signed(2, 8),
    to_signed(3, 8),
    to_signed(2, 8),
    to_signed(2, 8),
    to_signed(1, 8),
    to_signed(1, 8),
    to_signed(1, 8),
    to_signed(0, 8),
    to_signed(-2, 8),
    to_signed(-4, 8),
    to_signed(-6, 8),
    to_signed(-7, 8),
    to_signed(-7, 8),
    to_signed(-5, 8),
    to_signed(-2, 8),
    to_signed(0, 8),
    to_signed(1, 8),
    to_signed(2, 8),
    to_signed(1, 8),
    to_signed(0, 8),
    to_signed(-1, 8),
    to_signed(-2, 8),
    to_signed(-3, 8),
    to_signed(-3, 8),
    to_signed(-2, 8),
    to_signed(-1, 8),
    to_signed(0, 8),
    to_signed(0, 8),
    to_signed(0, 8),
    to_signed(-1, 8),
    to_signed(-2, 8),
    to_signed(-4, 8),
    to_signed(-6, 8),
    to_signed(-6, 8),
    to_signed(-5, 8),
    to_signed(-3, 8),
    to_signed(-2, 8),
    to_signed(-1, 8),
    to_signed(-1, 8),
    to_signed(-1, 8),
    to_signed(-2, 8),
    to_signed(-3, 8),
    to_signed(-3, 8),
    to_signed(-3, 8),
    to_signed(-2, 8),
    to_signed(-1, 8),
    to_signed(-1, 8),
    to_signed(0, 8),
    to_signed(1, 8),
    to_signed(2, 8),
    to_signed(1, 8),
    to_signed(0, 8),
    to_signed(-1, 8),
    to_signed(-2, 8),
    to_signed(-3, 8),
    to_signed(-2, 8),
    to_signed(-1, 8),
    to_signed(1, 8),
    to_signed(2, 8),
    to_signed(3, 8),
    to_signed(4, 8),
    to_signed(4, 8),
    to_signed(3, 8),
    to_signed(2, 8),
    to_signed(0, 8),
    to_signed(0, 8),
    to_signed(0, 8),
    to_signed(1, 8),
    to_signed(2, 8),
    to_signed(3, 8),
    to_signed(3, 8),
    to_signed(3, 8),
    to_signed(2, 8),
    to_signed(-1, 8),
    to_signed(-5, 8),
    to_signed(-9, 8),
    to_signed(-10, 8),
    to_signed(-8, 8),
    to_signed(-6, 8),
    to_signed(-4, 8),
    to_signed(-2, 8),
    to_signed(-1, 8),
    to_signed(-1, 8),
    to_signed(-2, 8),
    to_signed(-3, 8),
    to_signed(-5, 8),
    to_signed(-5, 8),
    to_signed(-4, 8),
    to_signed(-3, 8),
    to_signed(-1, 8),
    to_signed(0, 8),
    to_signed(0, 8),
    to_signed(0, 8),
    to_signed(0, 8),
    to_signed(-1, 8),
    to_signed(-2, 8),
    to_signed(-3, 8),
    to_signed(-4, 8),
    to_signed(-4, 8),
    to_signed(-3, 8),
    to_signed(-1, 8),
    to_signed(1, 8),
    to_signed(2, 8),
    to_signed(3, 8),
    to_signed(4, 8),
    to_signed(3, 8),
    to_signed(2, 8),
    to_signed(2, 8),
    to_signed(2, 8),
    to_signed(2, 8),
    to_signed(3, 8),
    to_signed(3, 8),
    to_signed(4, 8),
    to_signed(4, 8),
    to_signed(4, 8),
    to_signed(4, 8),
    to_signed(3, 8),
    to_signed(2, 8),
    to_signed(-1, 8),
    to_signed(-4, 8),
    to_signed(-6, 8),
    to_signed(-6, 8),
    to_signed(-5, 8),
    to_signed(-2, 8),
    to_signed(0, 8),
    to_signed(2, 8),
    to_signed(2, 8),
    to_signed(2, 8),
    to_signed(0, 8),
    to_signed(-1, 8),
    to_signed(-2, 8),
    to_signed(-2, 8),
    to_signed(-1, 8),
    to_signed(1, 8),
    to_signed(2, 8),
    to_signed(3, 8),
    to_signed(3, 8),
    to_signed(2, 8),
    to_signed(1, 8),
    to_signed(0, 8),
    to_signed(-1, 8),
    to_signed(-1, 8),
    to_signed(-2, 8),
    to_signed(-2, 8),
    to_signed(-2, 8),
    to_signed(-1, 8),
    to_signed(-1, 8),
    to_signed(0, 8),
    to_signed(1, 8),
    to_signed(2, 8),
    to_signed(3, 8),
    to_signed(3, 8),
    to_signed(3, 8),
    to_signed(3, 8),
    to_signed(2, 8),
    to_signed(2, 8),
    to_signed(2, 8),
    to_signed(4, 8),
    to_signed(5, 8),
    to_signed(6, 8),
    to_signed(6, 8),
    to_signed(6, 8),
    to_signed(4, 8),
    to_signed(3, 8),
    to_signed(1, 8),
    to_signed(1, 8),
    to_signed(2, 8),
    to_signed(3, 8),
    to_signed(4, 8),
    to_signed(6, 8),
    to_signed(7, 8),
    to_signed(7, 8),
    to_signed(8, 8),
    to_signed(7, 8),
    to_signed(7, 8),
    to_signed(7, 8),
    to_signed(7, 8),
    to_signed(7, 8),
    to_signed(6, 8),
    to_signed(6, 8),
    to_signed(6, 8),
    to_signed(6, 8),
    to_signed(6, 8),
    to_signed(4, 8),
    to_signed(2, 8),
    to_signed(0, 8),
    to_signed(-3, 8),
    to_signed(-3, 8),
    to_signed(-3, 8),
    to_signed(-1, 8),
    to_signed(1, 8),
    to_signed(3, 8),
    to_signed(3, 8),
    to_signed(2, 8),
    to_signed(1, 8),
    to_signed(0, 8),
    to_signed(0, 8),
    to_signed(0, 8),
    to_signed(2, 8),
    to_signed(3, 8),
    to_signed(4, 8),
    to_signed(4, 8),
    to_signed(4, 8),
    to_signed(4, 8),
    to_signed(4, 8),
    to_signed(3, 8),
    to_signed(1, 8),
    to_signed(-1, 8),
    to_signed(-2, 8),
    to_signed(-2, 8),
    to_signed(-1, 8),
    to_signed(1, 8),
    to_signed(3, 8),
    to_signed(4, 8),
    to_signed(6, 8),
    to_signed(7, 8),
    to_signed(8, 8),
    to_signed(7, 8),
    to_signed(7, 8),
    to_signed(8, 8),
    to_signed(9, 8),
    to_signed(9, 8),
    to_signed(9, 8),
    to_signed(10, 8),
    to_signed(10, 8),
    to_signed(9, 8),
    to_signed(8, 8),
    to_signed(7, 8),
    to_signed(6, 8),
    to_signed(4, 8),
    to_signed(3, 8),
    to_signed(3, 8),
    to_signed(3, 8),
    to_signed(4, 8),
    to_signed(4, 8),
    to_signed(5, 8),
    to_signed(4, 8),
    to_signed(3, 8),
    to_signed(2, 8),
    to_signed(0, 8),
    to_signed(-1, 8),
    to_signed(-2, 8),
    to_signed(-1, 8),
    to_signed(0, 8),
    to_signed(0, 8),
    to_signed(1, 8),
    to_signed(1, 8),
    to_signed(0, 8),
    to_signed(-2, 8),
    to_signed(-4, 8),
    to_signed(-6, 8),
    to_signed(-7, 8),
    to_signed(-7, 8),
    to_signed(-6, 8),
    to_signed(-4, 8),
    to_signed(-2, 8),
    to_signed(0, 8),
    to_signed(1, 8),
    to_signed(0, 8),
    to_signed(0, 8),
    to_signed(0, 8),
    to_signed(0, 8),
    to_signed(1, 8),
    to_signed(3, 8),
    to_signed(5, 8),
    to_signed(6, 8),
    to_signed(6, 8),
    to_signed(6, 8),
    to_signed(6, 8),
    to_signed(6, 8),
    to_signed(5, 8),
    to_signed(4, 8),
    to_signed(3, 8),
    to_signed(2, 8),
    to_signed(2, 8),
    to_signed(3, 8),
    to_signed(4, 8),
    to_signed(6, 8),
    to_signed(7, 8),
    to_signed(7, 8),
    to_signed(7, 8),
    to_signed(6, 8),
    to_signed(6, 8),
    to_signed(5, 8),
    to_signed(5, 8),
    to_signed(6, 8),
    to_signed(7, 8),
    to_signed(7, 8),
    to_signed(8, 8),
    to_signed(8, 8),
    to_signed(8, 8),
    to_signed(7, 8),
    to_signed(6, 8),
    to_signed(4, 8),
    to_signed(1, 8),
    to_signed(-1, 8),
    to_signed(-3, 8),
    to_signed(-3, 8),
    to_signed(-2, 8),
    to_signed(-1, 8),
    to_signed(0, 8),
    to_signed(0, 8),
    to_signed(-1, 8),
    to_signed(-2, 8),
    to_signed(-3, 8),
    to_signed(-4, 8),
    to_signed(-5, 8),
    to_signed(-5, 8),
    to_signed(-3, 8),
    to_signed(-2, 8),
    to_signed(-2, 8),
    to_signed(-2, 8),
    to_signed(-2, 8),
    to_signed(-3, 8),
    to_signed(-3, 8),
    to_signed(-4, 8),
    to_signed(-5, 8),
    to_signed(-6, 8),
    to_signed(-6, 8),
    to_signed(-6, 8),
    to_signed(-5, 8),
    to_signed(-5, 8),
    to_signed(-4, 8),
    to_signed(-3, 8),
    to_signed(-2, 8),
    to_signed(-1, 8),
    to_signed(-1, 8),
    to_signed(-1, 8),
    to_signed(-1, 8),
    to_signed(0, 8),
    to_signed(1, 8),
    to_signed(2, 8),
    to_signed(2, 8),
    to_signed(2, 8),
    to_signed(2, 8),
    to_signed(2, 8),
    to_signed(2, 8),
    to_signed(1, 8),
    to_signed(0, 8),
    to_signed(-2, 8),
    to_signed(-4, 8),
    to_signed(-4, 8),
    to_signed(-4, 8),
    to_signed(-4, 8),
    to_signed(-4, 8),
    to_signed(-4, 8),
    to_signed(-4, 8),
    to_signed(-4, 8),
    to_signed(-5, 8),
    to_signed(-5, 8),
    to_signed(-6, 8),
    to_signed(-6, 8),
    to_signed(-6, 8),
    to_signed(-5, 8),
    to_signed(-5, 8),
    to_signed(-6, 8),
    to_signed(-7, 8),
    to_signed(-8, 8),
    to_signed(-8, 8),
    to_signed(-9, 8),
    to_signed(-10, 8),
    to_signed(-11, 8),
    to_signed(-12, 8),
    to_signed(-12, 8),
    to_signed(-12, 8),
    to_signed(-11, 8),
    to_signed(-10, 8),
    to_signed(-9, 8),
    to_signed(-9, 8),
    to_signed(-9, 8),
    to_signed(-9, 8),
    to_signed(-8, 8),
    to_signed(-7, 8),
    to_signed(-5, 8),
    to_signed(-3, 8),
    to_signed(-2, 8),
    to_signed(-2, 8),
    to_signed(-3, 8),
    to_signed(-3, 8),
    to_signed(-3, 8),
    to_signed(-3, 8),
    to_signed(-3, 8),
    to_signed(-3, 8),
    to_signed(-4, 8),
    to_signed(-4, 8),
    to_signed(-3, 8),
    to_signed(-3, 8),
    to_signed(-3, 8),
    to_signed(-2, 8),
    to_signed(-2, 8),
    to_signed(-1, 8),
    to_signed(-1, 8),
    to_signed(-1, 8),
    to_signed(-1, 8),
    to_signed(-1, 8),
    to_signed(-1, 8),
    to_signed(0, 8),
    to_signed(0, 8),
    to_signed(0, 8),
    to_signed(0, 8),
    to_signed(0, 8),
    to_signed(0, 8),
    to_signed(-1, 8),
    to_signed(-2, 8),
    to_signed(-2, 8),
    to_signed(-3, 8),
    to_signed(-3, 8),
    to_signed(-3, 8),
    to_signed(-3, 8),
    to_signed(-3, 8),
    to_signed(-2, 8),
    to_signed(-2, 8),
    to_signed(-1, 8),
    to_signed(-1, 8),
    to_signed(0, 8),
    to_signed(1, 8),
    to_signed(1, 8),
    to_signed(1, 8),
    to_signed(2, 8),
    to_signed(2, 8),
    to_signed(1, 8),
    to_signed(0, 8),
    to_signed(0, 8),
    to_signed(-1, 8),
    to_signed(-2, 8),
    to_signed(-2, 8),
    to_signed(-3, 8),
    to_signed(-4, 8),
    to_signed(-5, 8),
    to_signed(-6, 8),
    to_signed(-6, 8),
    to_signed(-6, 8),
    to_signed(-6, 8),
    to_signed(-6, 8),
    to_signed(-6, 8),
    to_signed(-6, 8),
    to_signed(-4, 8),
    to_signed(-3, 8),
    to_signed(-1, 8),
    to_signed(0, 8),
    to_signed(1, 8),
    to_signed(1, 8),
    to_signed(1, 8),
    to_signed(0, 8),
    to_signed(0, 8),
    to_signed(0, 8),
    to_signed(0, 8),
    to_signed(0, 8),
    to_signed(0, 8),
    to_signed(0, 8),
    to_signed(0, 8),
    to_signed(-1, 8),
    to_signed(-1, 8),
    to_signed(-1, 8),
    to_signed(0, 8),
    to_signed(0, 8),
    to_signed(-1, 8),
    to_signed(-1, 8),
    to_signed(-2, 8),
    to_signed(-1, 8),
    to_signed(-1, 8),
    to_signed(0, 8),
    to_signed(1, 8),
    to_signed(0, 8),
    to_signed(0, 8),
    to_signed(-1, 8),
    to_signed(-3, 8),
    to_signed(-4, 8),
    to_signed(-5, 8),
    to_signed(-5, 8),
    to_signed(-5, 8),
    to_signed(-6, 8),
    to_signed(-7, 8),
    to_signed(-8, 8),
    to_signed(-10, 8),
    to_signed(-10, 8),
    to_signed(-10, 8),
    to_signed(-10, 8),
    to_signed(-9, 8),
    to_signed(-9, 8),
    to_signed(-8, 8),
    to_signed(-7, 8),
    to_signed(-7, 8),
    to_signed(-7, 8),
    to_signed(-5, 8),
    to_signed(-4, 8),
    to_signed(-4, 8),
    to_signed(-4, 8),
    to_signed(-5, 8),
    to_signed(-5, 8),
    to_signed(-5, 8),
    to_signed(-4, 8),
    to_signed(-3, 8),
    to_signed(-3, 8),
    to_signed(-2, 8),
    to_signed(-2, 8),
    to_signed(-3, 8),
    to_signed(-3, 8),
    to_signed(-4, 8),
    to_signed(-4, 8),
    to_signed(-4, 8),
    to_signed(-3, 8),
    to_signed(-1, 8),
    to_signed(1, 8),
    to_signed(3, 8),
    to_signed(4, 8),
    to_signed(5, 8),
    to_signed(4, 8),
    to_signed(4, 8),
    to_signed(3, 8),
    to_signed(2, 8),
    to_signed(1, 8),
    to_signed(0, 8),
    to_signed(0, 8),
    to_signed(-1, 8),
    to_signed(-1, 8),
    to_signed(-2, 8),
    to_signed(-3, 8),
    to_signed(-4, 8),
    to_signed(-4, 8),
    to_signed(-5, 8),
    to_signed(-5, 8),
    to_signed(-6, 8),
    to_signed(-6, 8),
    to_signed(-5, 8),
    to_signed(-4, 8),
    to_signed(-3, 8),
    to_signed(-2, 8),
    to_signed(-1, 8),
    to_signed(-2, 8),
    to_signed(-2, 8),
    to_signed(-3, 8),
    to_signed(-3, 8),
    to_signed(-3, 8),
    to_signed(-4, 8),
    to_signed(-3, 8),
    to_signed(-3, 8),
    to_signed(-2, 8),
    to_signed(-3, 8),
    to_signed(-3, 8),
    to_signed(-4, 8),
    to_signed(-4, 8),
    to_signed(-4, 8),
    to_signed(-4, 8),
    to_signed(-4, 8),
    to_signed(-4, 8),
    to_signed(-3, 8),
    to_signed(-1, 8),
    to_signed(0, 8),
    to_signed(2, 8),
    to_signed(3, 8),
    to_signed(3, 8),
    to_signed(2, 8),
    to_signed(1, 8),
    to_signed(0, 8),
    to_signed(-1, 8),
    to_signed(-1, 8),
    to_signed(0, 8),
    to_signed(1, 8),
    to_signed(1, 8),
    to_signed(1, 8),
    to_signed(0, 8),
    to_signed(-2, 8),
    to_signed(-3, 8),
    to_signed(-4, 8),
    to_signed(-5, 8),
    to_signed(-6, 8),
    to_signed(-6, 8),
    to_signed(-6, 8),
    to_signed(-5, 8),
    to_signed(-4, 8),
    to_signed(-3, 8),
    to_signed(-2, 8),
    to_signed(-1, 8),
    to_signed(0, 8),
    to_signed(-1, 8),
    to_signed(-1, 8),
    to_signed(-3, 8),
    to_signed(-4, 8),
    to_signed(-4, 8),
    to_signed(-3, 8),
    to_signed(-2, 8),
    to_signed(-1, 8),
    to_signed(-2, 8),
    to_signed(-2, 8),
    to_signed(-3, 8),
    to_signed(-4, 8),
    to_signed(-4, 8),
    to_signed(-5, 8),
    to_signed(-5, 8),
    to_signed(-4, 8),
    to_signed(-3, 8),
    to_signed(-1, 8),
    to_signed(1, 8),
    to_signed(2, 8),
    to_signed(3, 8),
    to_signed(3, 8),
    to_signed(3, 8),
    to_signed(2, 8),
    to_signed(1, 8),
    to_signed(0, 8),
    to_signed(0, 8),
    to_signed(1, 8),
    to_signed(2, 8),
    to_signed(2, 8),
    to_signed(1, 8),
    to_signed(0, 8),
    to_signed(-1, 8),
    to_signed(-2, 8),
    to_signed(-3, 8),
    to_signed(-4, 8),
    to_signed(-4, 8),
    to_signed(-3, 8),
    to_signed(-2, 8),
    to_signed(-1, 8),
    to_signed(1, 8),
    to_signed(2, 8),
    to_signed(2, 8),
    to_signed(1, 8),
    to_signed(1, 8),
    to_signed(0, 8),
    to_signed(-1, 8),
    to_signed(-1, 8),
    to_signed(-1, 8),
    to_signed(-1, 8),
    to_signed(-1, 8),
    to_signed(-2, 8),
    to_signed(-2, 8),
    to_signed(-3, 8),
    to_signed(-3, 8),
    to_signed(-4, 8),
    to_signed(-4, 8),
    to_signed(-5, 8),
    to_signed(-6, 8),
    to_signed(-6, 8),
    to_signed(-4, 8),
    to_signed(-3, 8),
    to_signed(-1, 8),
    to_signed(0, 8),
    to_signed(0, 8),
    to_signed(0, 8),
    to_signed(0, 8),
    to_signed(-1, 8),
    to_signed(-2, 8),
    to_signed(-3, 8),
    to_signed(-3, 8),
    to_signed(-2, 8),
    to_signed(-2, 8),
    to_signed(-2, 8),
    to_signed(-2, 8),
    to_signed(-3, 8),
    to_signed(-3, 8),
    to_signed(-2, 8),
    to_signed(-2, 8),
    to_signed(-2, 8),
    to_signed(-2, 8),
    to_signed(-1, 8),
    to_signed(0, 8),
    to_signed(2, 8),
    to_signed(3, 8),
    to_signed(4, 8),
    to_signed(5, 8),
    to_signed(5, 8),
    to_signed(5, 8),
    to_signed(4, 8),
    to_signed(3, 8),
    to_signed(2, 8),
    to_signed(1, 8),
    to_signed(1, 8),
    to_signed(1, 8),
    to_signed(0, 8),
    to_signed(0, 8),
    to_signed(-1, 8),
    to_signed(-2, 8),
    to_signed(-3, 8),
    to_signed(-4, 8),
    to_signed(-5, 8),
    to_signed(-6, 8),
    to_signed(-6, 8),
    to_signed(-6, 8),
    to_signed(-5, 8),
    to_signed(-5, 8),
    to_signed(-4, 8),
    to_signed(-3, 8),
    to_signed(-3, 8),
    to_signed(-3, 8),
    to_signed(-4, 8),
    to_signed(-5, 8),
    to_signed(-7, 8),
    to_signed(-8, 8),
    to_signed(-9, 8),
    to_signed(-9, 8),
    to_signed(-9, 8),
    to_signed(-9, 8),
    to_signed(-9, 8),
    to_signed(-9, 8),
    to_signed(-10, 8),
    to_signed(-10, 8),
    to_signed(-10, 8),
    to_signed(-10, 8),
    to_signed(-10, 8),
    to_signed(-8, 8),
    to_signed(-7, 8),
    to_signed(-5, 8),
    to_signed(-4, 8),
    to_signed(-3, 8),
    to_signed(-2, 8),
    to_signed(-1, 8),
    to_signed(0, 8),
    to_signed(0, 8),
    to_signed(1, 8),
    to_signed(1, 8),
    to_signed(1, 8),
    to_signed(1, 8),
    to_signed(1, 8),
    to_signed(1, 8),
    to_signed(0, 8),
    to_signed(0, 8),
    to_signed(0, 8),
    to_signed(-1, 8),
    to_signed(-2, 8),
    to_signed(-3, 8),
    to_signed(-3, 8),
    to_signed(-3, 8),
    to_signed(-2, 8),
    to_signed(-2, 8),
    to_signed(-2, 8),
    to_signed(-2, 8),
    to_signed(-2, 8),
    to_signed(-2, 8),
    to_signed(-2, 8),
    to_signed(-3, 8),
    to_signed(-4, 8),
    to_signed(-5, 8),
    to_signed(-5, 8),
    to_signed(-5, 8),
    to_signed(-5, 8),
    to_signed(-5, 8),
    to_signed(-5, 8),
    to_signed(-5, 8),
    to_signed(-5, 8),
    to_signed(-5, 8),
    to_signed(-5, 8),
    to_signed(-6, 8),
    to_signed(-5, 8),
    to_signed(-5, 8),
    to_signed(-3, 8),
    to_signed(-2, 8),
    to_signed(-2, 8),
    to_signed(0, 8),
    to_signed(1, 8),
    to_signed(2, 8),
    to_signed(3, 8),
    to_signed(3, 8),
    to_signed(2, 8),
    to_signed(2, 8),
    to_signed(3, 8),
    to_signed(3, 8),
    to_signed(3, 8),
    to_signed(4, 8),
    to_signed(4, 8),
    to_signed(5, 8),
    to_signed(5, 8),
    to_signed(6, 8),
    to_signed(6, 8),
    to_signed(6, 8),
    to_signed(7, 8),
    to_signed(8, 8),
    to_signed(9, 8),
    to_signed(10, 8),
    to_signed(10, 8),
    to_signed(11, 8),
    to_signed(12, 8),
    to_signed(13, 8),
    to_signed(14, 8),
    to_signed(14, 8),
    to_signed(13, 8),
    to_signed(12, 8),
    to_signed(11, 8),
    to_signed(10, 8),
    to_signed(9, 8),
    to_signed(8, 8),
    to_signed(7, 8),
    to_signed(7, 8),
    to_signed(6, 8),
    to_signed(5, 8),
    to_signed(4, 8),
    to_signed(4, 8),
    to_signed(4, 8),
    to_signed(4, 8),
    to_signed(4, 8),
    to_signed(4, 8),
    to_signed(5, 8),
    to_signed(5, 8),
    to_signed(6, 8),
    to_signed(6, 8),
    to_signed(6, 8),
    to_signed(5, 8),
    to_signed(4, 8),
    to_signed(3, 8),
    to_signed(3, 8),
    to_signed(3, 8),
    to_signed(2, 8),
    to_signed(1, 8),
    to_signed(1, 8),
    to_signed(1, 8),
    to_signed(1, 8),
    to_signed(0, 8),
    to_signed(0, 8),
    to_signed(1, 8),
    to_signed(2, 8),
    to_signed(3, 8),
    to_signed(4, 8),
    to_signed(4, 8),
    to_signed(4, 8),
    to_signed(5, 8),
    to_signed(6, 8),
    to_signed(7, 8),
    to_signed(8, 8),
    to_signed(9, 8),
    to_signed(9, 8),
    to_signed(9, 8),
    to_signed(9, 8),
    to_signed(9, 8),
    to_signed(9, 8),
    to_signed(9, 8),
    to_signed(9, 8),
    to_signed(9, 8),
    to_signed(9, 8),
    to_signed(9, 8),
    to_signed(9, 8),
    to_signed(9, 8),
    to_signed(9, 8),
    to_signed(9, 8),
    to_signed(8, 8),
    to_signed(8, 8),
    to_signed(7, 8),
    to_signed(7, 8),
    to_signed(8, 8),
    to_signed(9, 8),
    to_signed(9, 8),
    to_signed(8, 8),
    to_signed(7, 8),
    to_signed(6, 8),
    to_signed(5, 8),
    to_signed(4, 8),
    to_signed(3, 8),
    to_signed(2, 8),
    to_signed(2, 8),
    to_signed(1, 8),
    to_signed(-1, 8),
    to_signed(-2, 8),
    to_signed(-2, 8),
    to_signed(-2, 8),
    to_signed(-2, 8),
    to_signed(-2, 8),
    to_signed(-2, 8),
    to_signed(-2, 8),
    to_signed(-2, 8),
    to_signed(-1, 8),
    to_signed(0, 8),
    to_signed(1, 8),
    to_signed(1, 8),
    to_signed(2, 8),
    to_signed(2, 8),
    to_signed(2, 8),
    to_signed(2, 8),
    to_signed(2, 8),
    to_signed(2, 8),
    to_signed(2, 8),
    to_signed(3, 8),
    to_signed(3, 8),
    to_signed(3, 8),
    to_signed(3, 8),
    to_signed(3, 8),
    to_signed(4, 8),
    to_signed(5, 8),
    to_signed(5, 8),
    to_signed(6, 8),
    to_signed(6, 8),
    to_signed(6, 8),
    to_signed(7, 8),
    to_signed(8, 8),
    to_signed(8, 8),
    to_signed(8, 8),
    to_signed(8, 8),
    to_signed(8, 8),
    to_signed(8, 8),
    to_signed(7, 8),
    to_signed(7, 8),
    to_signed(6, 8),
    to_signed(5, 8),
    to_signed(5, 8),
    to_signed(4, 8),
    to_signed(2, 8),
    to_signed(1, 8),
    to_signed(1, 8),
    to_signed(1, 8),
    to_signed(1, 8),
    to_signed(0, 8),
    to_signed(-1, 8),
    to_signed(-1, 8),
    to_signed(-2, 8),
    to_signed(-2, 8),
    to_signed(-1, 8),
    to_signed(-1, 8),
    to_signed(-1, 8),
    to_signed(-2, 8),
    to_signed(-3, 8),
    to_signed(-4, 8),
    to_signed(-5, 8),
    to_signed(-5, 8),
    to_signed(-6, 8),
    to_signed(-6, 8),
    to_signed(-6, 8),
    to_signed(-6, 8),
    to_signed(-7, 8),
    to_signed(-8, 8),
    to_signed(-8, 8),
    to_signed(-8, 8),
    to_signed(-9, 8),
    to_signed(-9, 8),
    to_signed(-8, 8),
    to_signed(-7, 8),
    to_signed(-7, 8),
    to_signed(-6, 8),
    to_signed(-4, 8),
    to_signed(-3, 8),
    to_signed(-2, 8),
    to_signed(-2, 8),
    to_signed(-1, 8),
    to_signed(-1, 8),
    to_signed(-1, 8),
    to_signed(-1, 8),
    to_signed(-1, 8),
    to_signed(-1, 8),
    to_signed(0, 8),
    to_signed(0, 8),
    to_signed(1, 8),
    to_signed(1, 8),
    to_signed(1, 8),
    to_signed(1, 8),
    to_signed(1, 8),
    to_signed(0, 8),
    to_signed(-1, 8),
    to_signed(-1, 8),
    to_signed(-2, 8),
    to_signed(-1, 8),
    to_signed(0, 8),
    to_signed(0, 8),
    to_signed(0, 8),
    to_signed(0, 8),
    to_signed(-1, 8),
    to_signed(-2, 8),
    to_signed(-3, 8),
    to_signed(-4, 8),
    to_signed(-6, 8),
    to_signed(-7, 8),
    to_signed(-8, 8),
    to_signed(-9, 8),
    to_signed(-10, 8),
    to_signed(-10, 8),
    to_signed(-10, 8),
    to_signed(-10, 8),
    to_signed(-10, 8),
    to_signed(-11, 8),
    to_signed(-12, 8),
    to_signed(-13, 8),
    to_signed(-13, 8),
    to_signed(-12, 8),
    to_signed(-11, 8),
    to_signed(-9, 8),
    to_signed(-8, 8),
    to_signed(-7, 8),
    to_signed(-7, 8),
    to_signed(-7, 8),
    to_signed(-7, 8),
    to_signed(-7, 8),
    to_signed(-7, 8),
    to_signed(-6, 8),
    to_signed(-6, 8),
    to_signed(-4, 8),
    to_signed(-4, 8),
    to_signed(-3, 8),
    to_signed(-1, 8),
    to_signed(-1, 8),
    to_signed(0, 8),
    to_signed(0, 8),
    to_signed(0, 8),
    to_signed(1, 8),
    to_signed(1, 8),
    to_signed(3, 8),
    to_signed(4, 8),
    to_signed(5, 8),
    to_signed(6, 8),
    to_signed(7, 8),
    to_signed(7, 8),
    to_signed(6, 8),
    to_signed(6, 8),
    to_signed(5, 8),
    to_signed(4, 8),
    to_signed(3, 8),
    to_signed(2, 8),
    to_signed(1, 8),
    to_signed(1, 8),
    to_signed(0, 8),
    to_signed(0, 8),
    to_signed(0, 8),
    to_signed(-1, 8),
    to_signed(-2, 8),
    to_signed(-4, 8),
    to_signed(-5, 8),
    to_signed(-6, 8),
    to_signed(-6, 8),
    to_signed(-6, 8),
    to_signed(-5, 8),
    to_signed(-4, 8),
    to_signed(-4, 8),
    to_signed(-4, 8),
    to_signed(-5, 8),
    to_signed(-6, 8),
    to_signed(-6, 8),
    to_signed(-7, 8),
    to_signed(-7, 8),
    to_signed(-7, 8),
    to_signed(-7, 8),
    to_signed(-7, 8),
    to_signed(-7, 8),
    to_signed(-7, 8),
    to_signed(-7, 8),
    to_signed(-6, 8),
    to_signed(-5, 8),
    to_signed(-3, 8),
    to_signed(-2, 8),
    to_signed(-1, 8),
    to_signed(0, 8),
    to_signed(2, 8),
    to_signed(4, 8),
    to_signed(5, 8),
    to_signed(7, 8),
    to_signed(8, 8),
    to_signed(10, 8),
    to_signed(11, 8),
    to_signed(11, 8),
    to_signed(10, 8),
    to_signed(9, 8),
    to_signed(8, 8),
    to_signed(8, 8),
    to_signed(8, 8),
    to_signed(8, 8),
    to_signed(9, 8),
    to_signed(9, 8),
    to_signed(9, 8),
    to_signed(9, 8),
    to_signed(8, 8),
    to_signed(6, 8),
    to_signed(5, 8),
    to_signed(5, 8),
    to_signed(6, 8),
    to_signed(7, 8),
    to_signed(7, 8),
    to_signed(7, 8),
    to_signed(6, 8),
    to_signed(5, 8),
    to_signed(5, 8),
    to_signed(3, 8),
    to_signed(2, 8),
    to_signed(0, 8),
    to_signed(-1, 8),
    to_signed(-2, 8),
    to_signed(-3, 8),
    to_signed(-4, 8),
    to_signed(-4, 8),
    to_signed(-5, 8),
    to_signed(-5, 8),
    to_signed(-6, 8),
    to_signed(-8, 8),
    to_signed(-9, 8),
    to_signed(-10, 8),
    to_signed(-9, 8),
    to_signed(-7, 8),
    to_signed(-5, 8),
    to_signed(-4, 8),
    to_signed(-4, 8),
    to_signed(-3, 8),
    to_signed(-3, 8),
    to_signed(-3, 8),
    to_signed(-3, 8),
    to_signed(-3, 8),
    to_signed(-2, 8),
    to_signed(-1, 8),
    to_signed(-1, 8),
    to_signed(-1, 8),
    to_signed(0, 8),
    to_signed(0, 8),
    to_signed(1, 8),
    to_signed(2, 8),
    to_signed(2, 8),
    to_signed(2, 8),
    to_signed(3, 8),
    to_signed(4, 8),
    to_signed(5, 8),
    to_signed(7, 8),
    to_signed(9, 8),
    to_signed(10, 8),
    to_signed(11, 8),
    to_signed(11, 8),
    to_signed(12, 8),
    to_signed(12, 8),
    to_signed(11, 8),
    to_signed(10, 8),
    to_signed(9, 8),
    to_signed(8, 8),
    to_signed(7, 8),
    to_signed(6, 8),
    to_signed(6, 8),
    to_signed(6, 8),
    to_signed(5, 8),
    to_signed(5, 8),
    to_signed(4, 8),
    to_signed(3, 8),
    to_signed(2, 8),
    to_signed(0, 8),
    to_signed(0, 8),
    to_signed(0, 8),
    to_signed(0, 8),
    to_signed(1, 8),
    to_signed(1, 8),
    to_signed(1, 8),
    to_signed(1, 8),
    to_signed(0, 8),
    to_signed(-1, 8),
    to_signed(-2, 8),
    to_signed(-3, 8),
    to_signed(-4, 8),
    to_signed(-5, 8),
    to_signed(-5, 8),
    to_signed(-5, 8),
    to_signed(-5, 8),
    to_signed(-5, 8),
    to_signed(-5, 8),
    to_signed(-5, 8),
    to_signed(-5, 8),
    to_signed(-5, 8),
    to_signed(-5, 8),
    to_signed(-5, 8),
    to_signed(-4, 8),
    to_signed(-3, 8),
    to_signed(-1, 8),
    to_signed(1, 8),
    to_signed(2, 8),
    to_signed(3, 8),
    to_signed(4, 8),
    to_signed(4, 8),
    to_signed(4, 8),
    to_signed(3, 8),
    to_signed(3, 8),
    to_signed(3, 8),
    to_signed(3, 8),
    to_signed(3, 8),
    to_signed(4, 8),
    to_signed(4, 8),
    to_signed(4, 8),
    to_signed(3, 8),
    to_signed(3, 8),
    to_signed(2, 8),
    to_signed(1, 8),
    to_signed(1, 8),
    to_signed(2, 8),
    to_signed(3, 8),
    to_signed(3, 8),
    to_signed(3, 8),
    to_signed(4, 8),
    to_signed(4, 8),
    to_signed(4, 8),
    to_signed(2, 8),
    to_signed(0, 8),
    to_signed(-1, 8),
    to_signed(-2, 8),
    to_signed(-3, 8),
    to_signed(-4, 8),
    to_signed(-4, 8),
    to_signed(-4, 8),
    to_signed(-4, 8),
    to_signed(-5, 8),
    to_signed(-6, 8),
    to_signed(-7, 8),
    to_signed(-8, 8),
    to_signed(-9, 8),
    to_signed(-8, 8),
    to_signed(-8, 8),
    to_signed(-7, 8),
    to_signed(-7, 8),
    to_signed(-6, 8),
    to_signed(-5, 8),
    to_signed(-4, 8),
    to_signed(-5, 8),
    to_signed(-5, 8),
    to_signed(-6, 8),
    to_signed(-6, 8),
    to_signed(-7, 8),
    to_signed(-7, 8),
    to_signed(-7, 8),
    to_signed(-6, 8),
    to_signed(-5, 8),
    to_signed(-4, 8),
    to_signed(-3, 8),
    to_signed(-3, 8),
    to_signed(-3, 8),
    to_signed(-3, 8),
    to_signed(-2, 8),
    to_signed(-2, 8),
    to_signed(-1, 8),
    to_signed(0, 8),
    to_signed(2, 8),
    to_signed(3, 8),
    to_signed(4, 8),
    to_signed(5, 8),
    to_signed(4, 8),
    to_signed(3, 8),
    to_signed(2, 8),
    to_signed(2, 8),
    to_signed(1, 8),
    to_signed(0, 8),
    to_signed(0, 8),
    to_signed(-1, 8),
    to_signed(-1, 8),
    to_signed(-1, 8),
    to_signed(-1, 8),
    to_signed(-2, 8),
    to_signed(-3, 8),
    to_signed(-3, 8),
    to_signed(-4, 8),
    to_signed(-4, 8),
    to_signed(-4, 8),
    to_signed(-4, 8),
    to_signed(-4, 8),
    to_signed(-3, 8),
    to_signed(-3, 8),
    to_signed(-3, 8),
    to_signed(-3, 8),
    to_signed(-3, 8),
    to_signed(-4, 8),
    to_signed(-5, 8),
    to_signed(-6, 8),
    to_signed(-7, 8),
    to_signed(-8, 8),
    to_signed(-8, 8),
    to_signed(-8, 8),
    to_signed(-8, 8),
    to_signed(-8, 8),
    to_signed(-7, 8),
    to_signed(-7, 8),
    to_signed(-7, 8),
    to_signed(-6, 8),
    to_signed(-6, 8),
    to_signed(-6, 8),
    to_signed(-6, 8),
    to_signed(-5, 8),
    to_signed(-4, 8),
    to_signed(-3, 8),
    to_signed(-2, 8),
    to_signed(-1, 8),
    to_signed(-1, 8),
    to_signed(-1, 8),
    to_signed(-2, 8),
    to_signed(-2, 8),
    to_signed(-3, 8),
    to_signed(-3, 8),
    to_signed(-3, 8),
    to_signed(-3, 8),
    to_signed(-3, 8),
    to_signed(-3, 8),
    to_signed(-3, 8),
    to_signed(-3, 8),
    to_signed(-3, 8),
    to_signed(-3, 8),
    to_signed(-4, 8),
    to_signed(-4, 8),
    to_signed(-4, 8),
    to_signed(-3, 8),
    to_signed(-3, 8),
    to_signed(-2, 8),
    to_signed(-1, 8),
    to_signed(-2, 8),
    to_signed(-2, 8),
    to_signed(-3, 8),
    to_signed(-5, 8),
    to_signed(-6, 8),
    to_signed(-8, 8),
    to_signed(-8, 8),
    to_signed(-8, 8),
    to_signed(-9, 8),
    to_signed(-9, 8),
    to_signed(-9, 8),
    to_signed(-9, 8),
    to_signed(-8, 8),
    to_signed(-8, 8),
    to_signed(-8, 8),
    to_signed(-8, 8),
    to_signed(-8, 8),
    to_signed(-8, 8),
    to_signed(-6, 8),
    to_signed(-5, 8),
    to_signed(-3, 8),
    to_signed(-2, 8),
    to_signed(-2, 8),
    to_signed(-2, 8),
    to_signed(-3, 8),
    to_signed(-4, 8),
    to_signed(-4, 8),
    to_signed(-4, 8),
    to_signed(-5, 8),
    to_signed(-5, 8),
    to_signed(-6, 8),
    to_signed(-6, 8),
    to_signed(-6, 8),
    to_signed(-5, 8),
    to_signed(-5, 8),
    to_signed(-5, 8),
    to_signed(-5, 8),
    to_signed(-5, 8),
    to_signed(-5, 8),
    to_signed(-4, 8),
    to_signed(-4, 8),
    to_signed(-2, 8),
    to_signed(-1, 8),
    to_signed(-1, 8),
    to_signed(-1, 8),
    to_signed(-1, 8),
    to_signed(-1, 8),
    to_signed(-2, 8),
    to_signed(-3, 8),
    to_signed(-3, 8),
    to_signed(-4, 8),
    to_signed(-4, 8),
    to_signed(-5, 8),
    to_signed(-5, 8),
    to_signed(-4, 8),
    to_signed(-4, 8),
    to_signed(-4, 8),
    to_signed(-4, 8),
    to_signed(-3, 8),
    to_signed(-3, 8),
    to_signed(-2, 8),
    to_signed(-2, 8),
    to_signed(-2, 8),
    to_signed(-1, 8),
    to_signed(0, 8),
    to_signed(1, 8),
    to_signed(1, 8),
    to_signed(1, 8),
    to_signed(1, 8),
    to_signed(0, 8),
    to_signed(0, 8),
    to_signed(0, 8),
    to_signed(-1, 8),
    to_signed(-1, 8),
    to_signed(-2, 8),
    to_signed(-3, 8),
    to_signed(-2, 8),
    to_signed(-1, 8),
    to_signed(-1, 8),
    to_signed(-1, 8),
    to_signed(-1, 8),
    to_signed(-2, 8),
    to_signed(-3, 8),
    to_signed(-4, 8),
    to_signed(-3, 8),
    to_signed(-2, 8),
    to_signed(0, 8),
    to_signed(1, 8),
    to_signed(1, 8),
    to_signed(0, 8),
    to_signed(0, 8),
    to_signed(-1, 8),
    to_signed(-1, 8),
    to_signed(-1, 8),
    to_signed(-2, 8),
    to_signed(-2, 8),
    to_signed(-2, 8),
    to_signed(-3, 8),
    to_signed(-2, 8),
    to_signed(-2, 8),
    to_signed(-1, 8),
    to_signed(-1, 8),
    to_signed(-1, 8),
    to_signed(-1, 8),
    to_signed(-2, 8),
    to_signed(-2, 8),
    to_signed(-1, 8),
    to_signed(1, 8),
    to_signed(3, 8),
    to_signed(5, 8),
    to_signed(5, 8),
    to_signed(5, 8),
    to_signed(4, 8),
    to_signed(4, 8),
    to_signed(3, 8),
    to_signed(3, 8),
    to_signed(3, 8),
    to_signed(3, 8),
    to_signed(2, 8),
    to_signed(1, 8),
    to_signed(1, 8),
    to_signed(1, 8),
    to_signed(1, 8),
    to_signed(1, 8),
    to_signed(1, 8),
    to_signed(1, 8),
    to_signed(1, 8),
    to_signed(1, 8),
    to_signed(2, 8),
    to_signed(2, 8),
    to_signed(2, 8),
    to_signed(3, 8),
    to_signed(3, 8),
    to_signed(2, 8),
    to_signed(2, 8),
    to_signed(1, 8),
    to_signed(0, 8),
    to_signed(-1, 8),
    to_signed(-1, 8),
    to_signed(-3, 8),
    to_signed(-4, 8),
    to_signed(-5, 8),
    to_signed(-5, 8),
    to_signed(-5, 8),
    to_signed(-5, 8),
    to_signed(-5, 8),
    to_signed(-6, 8),
    to_signed(-7, 8),
    to_signed(-7, 8),
    to_signed(-6, 8),
    to_signed(-5, 8),
    to_signed(-4, 8),
    to_signed(-3, 8),
    to_signed(-3, 8),
    to_signed(-3, 8),
    to_signed(-3, 8),
    to_signed(-4, 8),
    to_signed(-4, 8),
    to_signed(-4, 8),
    to_signed(-3, 8),
    to_signed(-4, 8),
    to_signed(-4, 8),
    to_signed(-5, 8),
    to_signed(-4, 8),
    to_signed(-4, 8),
    to_signed(-3, 8),
    to_signed(-2, 8),
    to_signed(-1, 8),
    to_signed(-1, 8),
    to_signed(-1, 8),
    to_signed(-1, 8),
    to_signed(0, 8),
    to_signed(1, 8),
    to_signed(2, 8),
    to_signed(4, 8),
    to_signed(4, 8),
    to_signed(4, 8),
    to_signed(4, 8),
    to_signed(3, 8),
    to_signed(3, 8),
    to_signed(3, 8),
    to_signed(3, 8),
    to_signed(3, 8),
    to_signed(1, 8),
    to_signed(0, 8),
    to_signed(-1, 8),
    to_signed(0, 8),
    to_signed(0, 8),
    to_signed(1, 8),
    to_signed(1, 8),
    to_signed(1, 8),
    to_signed(0, 8),
    to_signed(0, 8),
    to_signed(0, 8),
    to_signed(1, 8),
    to_signed(2, 8),
    to_signed(2, 8),
    to_signed(2, 8),
    to_signed(2, 8),
    to_signed(2, 8),
    to_signed(1, 8),
    to_signed(1, 8),
    to_signed(0, 8),
    to_signed(0, 8),
    to_signed(-1, 8),
    to_signed(-2, 8),
    to_signed(-3, 8),
    to_signed(-4, 8),
    to_signed(-4, 8),
    to_signed(-3, 8),
    to_signed(-3, 8),
    to_signed(-2, 8),
    to_signed(-2, 8),
    to_signed(-2, 8),
    to_signed(-1, 8),
    to_signed(0, 8),
    to_signed(2, 8),
    to_signed(3, 8),
    to_signed(4, 8),
    to_signed(5, 8),
    to_signed(6, 8),
    to_signed(6, 8),
    to_signed(6, 8),
    to_signed(6, 8),
    to_signed(6, 8),
    to_signed(6, 8),
    to_signed(5, 8),
    to_signed(5, 8),
    to_signed(4, 8),
    to_signed(4, 8),
    to_signed(4, 8),
    to_signed(5, 8),
    to_signed(5, 8),
    to_signed(5, 8),
    to_signed(5, 8),
    to_signed(5, 8),
    to_signed(6, 8),
    to_signed(8, 8),
    to_signed(9, 8),
    to_signed(10, 8),
    to_signed(11, 8),
    to_signed(12, 8),
    to_signed(12, 8),
    to_signed(11, 8),
    to_signed(10, 8),
    to_signed(10, 8),
    to_signed(9, 8),
    to_signed(8, 8),
    to_signed(7, 8),
    to_signed(5, 8),
    to_signed(4, 8),
    to_signed(3, 8),
    to_signed(2, 8),
    to_signed(2, 8),
    to_signed(2, 8),
    to_signed(2, 8),
    to_signed(0, 8),
    to_signed(0, 8),
    to_signed(0, 8),
    to_signed(0, 8),
    to_signed(1, 8),
    to_signed(1, 8),
    to_signed(2, 8),
    to_signed(3, 8),
    to_signed(3, 8),
    to_signed(2, 8),
    to_signed(2, 8),
    to_signed(1, 8),
    to_signed(1, 8),
    to_signed(0, 8),
    to_signed(-1, 8),
    to_signed(-3, 8),
    to_signed(-4, 8),
    to_signed(-4, 8),
    to_signed(-4, 8),
    to_signed(-4, 8),
    to_signed(-3, 8),
    to_signed(-2, 8),
    to_signed(-2, 8),
    to_signed(-2, 8),
    to_signed(-2, 8),
    to_signed(-1, 8),
    to_signed(1, 8),
    to_signed(1, 8),
    to_signed(2, 8),
    to_signed(3, 8),
    to_signed(3, 8),
    to_signed(4, 8),
    to_signed(4, 8),
    to_signed(5, 8),
    to_signed(5, 8),
    to_signed(4, 8),
    to_signed(3, 8),
    to_signed(1, 8),
    to_signed(0, 8),
    to_signed(-1, 8),
    to_signed(-1, 8),
    to_signed(-1, 8),
    to_signed(-1, 8),
    to_signed(-1, 8),
    to_signed(-1, 8),
    to_signed(-1, 8),
    to_signed(-1, 8),
    to_signed(-1, 8),
    to_signed(0, 8),
    to_signed(0, 8),
    to_signed(1, 8),
    to_signed(1, 8),
    to_signed(1, 8),
    to_signed(0, 8),
    to_signed(0, 8),
    to_signed(0, 8),
    to_signed(-1, 8),
    to_signed(-2, 8),
    to_signed(-3, 8),
    to_signed(-5, 8),
    to_signed(-6, 8),
    to_signed(-6, 8),
    to_signed(-6, 8),
    to_signed(-6, 8),
    to_signed(-5, 8),
    to_signed(-5, 8),
    to_signed(-6, 8),
    to_signed(-6, 8),
    to_signed(-5, 8),
    to_signed(-5, 8),
    to_signed(-4, 8),
    to_signed(-3, 8),
    to_signed(-2, 8),
    to_signed(-1, 8),
    to_signed(-1, 8),
    to_signed(0, 8),
    to_signed(0, 8),
    to_signed(0, 8),
    to_signed(0, 8),
    to_signed(0, 8),
    to_signed(0, 8),
    to_signed(-1, 8),
    to_signed(-2, 8),
    to_signed(-3, 8),
    to_signed(-3, 8),
    to_signed(-3, 8),
    to_signed(-3, 8),
    to_signed(-3, 8),
    to_signed(-4, 8),
    to_signed(-4, 8),
    to_signed(-3, 8),
    to_signed(-3, 8),
    to_signed(-2, 8),
    to_signed(-1, 8),
    to_signed(-1, 8),
    to_signed(-1, 8),
    to_signed(-1, 8),
    to_signed(-2, 8),
    to_signed(-2, 8),
    to_signed(-2, 8),
    to_signed(-2, 8),
    to_signed(-2, 8),
    to_signed(-3, 8),
    to_signed(-4, 8),
    to_signed(-5, 8),
    to_signed(-5, 8),
    to_signed(-5, 8),
    to_signed(-5, 8),
    to_signed(-5, 8),
    to_signed(-5, 8),
    to_signed(-5, 8),
    to_signed(-4, 8),
    to_signed(-3, 8),
    to_signed(-2, 8),
    to_signed(-1, 8),
    to_signed(0, 8),
    to_signed(1, 8),
    to_signed(2, 8),
    to_signed(2, 8),
    to_signed(3, 8),
    to_signed(3, 8),
    to_signed(3, 8),
    to_signed(4, 8),
    to_signed(4, 8),
    to_signed(3, 8),
    to_signed(1, 8),
    to_signed(0, 8),
    to_signed(-1, 8),
    to_signed(-1, 8),
    to_signed(1, 8),
    to_signed(2, 8),
    to_signed(2, 8),
    to_signed(1, 8),
    to_signed(1, 8),
    to_signed(2, 8),
    to_signed(4, 8),
    to_signed(5, 8),
    to_signed(5, 8),
    to_signed(3, 8),
    to_signed(2, 8),
    to_signed(2, 8),
    to_signed(2, 8),
    to_signed(2, 8),
    to_signed(2, 8),
    to_signed(2, 8),
    to_signed(2, 8),
    to_signed(1, 8),
    to_signed(0, 8),
    to_signed(-2, 8),
    to_signed(-3, 8),
    to_signed(-3, 8),
    to_signed(-3, 8),
    to_signed(-2, 8),
    to_signed(-3, 8),
    to_signed(-4, 8),
    to_signed(-4, 8),
    to_signed(-3, 8),
    to_signed(-1, 8),
    to_signed(0, 8),
    to_signed(0, 8),
    to_signed(1, 8),
    to_signed(1, 8),
    to_signed(1, 8),
    to_signed(1, 8),
    to_signed(1, 8),
    to_signed(1, 8),
    to_signed(0, 8),
    to_signed(0, 8),
    to_signed(-1, 8),
    to_signed(-1, 8),
    to_signed(-1, 8),
    to_signed(0, 8),
    to_signed(0, 8),
    to_signed(0, 8),
    to_signed(0, 8),
    to_signed(-1, 8),
    to_signed(-1, 8),
    to_signed(0, 8),
    to_signed(1, 8),
    to_signed(1, 8),
    to_signed(2, 8),
    to_signed(3, 8),
    to_signed(4, 8),
    to_signed(5, 8),
    to_signed(4, 8),
    to_signed(3, 8),
    to_signed(2, 8),
    to_signed(3, 8),
    to_signed(3, 8),
    to_signed(2, 8),
    to_signed(1, 8),
    to_signed(-1, 8),
    to_signed(-1, 8),
    to_signed(-2, 8),
    to_signed(-2, 8),
    to_signed(-2, 8),
    to_signed(-3, 8),
    to_signed(-3, 8),
    to_signed(-4, 8),
    to_signed(-4, 8),
    to_signed(-3, 8),
    to_signed(-3, 8),
    to_signed(-2, 8),
    to_signed(-1, 8),
    to_signed(-2, 8),
    to_signed(-2, 8),
    to_signed(-2, 8),
    to_signed(-2, 8),
    to_signed(-2, 8),
    to_signed(-2, 8),
    to_signed(-2, 8),
    to_signed(-3, 8),
    to_signed(-4, 8),
    to_signed(-5, 8),
    to_signed(-6, 8),
    to_signed(-6, 8),
    to_signed(-6, 8),
    to_signed(-5, 8),
    to_signed(-5, 8),
    to_signed(-6, 8),
    to_signed(-6, 8),
    to_signed(-5, 8),
    to_signed(-4, 8),
    to_signed(-3, 8),
    to_signed(-2, 8),
    to_signed(-2, 8),
    to_signed(-1, 8),
    to_signed(-1, 8),
    to_signed(-1, 8),
    to_signed(-1, 8),
    to_signed(-1, 8),
    to_signed(0, 8),
    to_signed(0, 8),
    to_signed(-1, 8),
    to_signed(-2, 8),
    to_signed(-3, 8),
    to_signed(-3, 8),
    to_signed(-3, 8),
    to_signed(-3, 8),
    to_signed(-3, 8),
    to_signed(-4, 8),
    to_signed(-4, 8),
    to_signed(-4, 8),
    to_signed(-4, 8),
    to_signed(-2, 8),
    to_signed(-1, 8),
    to_signed(-1, 8),
    to_signed(0, 8),
    to_signed(0, 8),
    to_signed(0, 8),
    to_signed(0, 8),
    to_signed(-1, 8),
    to_signed(-1, 8),
    to_signed(-1, 8),
    to_signed(-1, 8),
    to_signed(-1, 8),
    to_signed(-2, 8),
    to_signed(-2, 8),
    to_signed(-2, 8),
    to_signed(-2, 8),
    to_signed(-2, 8),
    to_signed(-2, 8),
    to_signed(-2, 8),
    to_signed(-2, 8),
    to_signed(-2, 8),
    to_signed(-2, 8),
    to_signed(-1, 8),
    to_signed(1, 8),
    to_signed(3, 8),
    to_signed(3, 8),
    to_signed(3, 8),
    to_signed(3, 8),
    to_signed(3, 8),
    to_signed(3, 8),
    to_signed(3, 8),
    to_signed(4, 8),
    to_signed(4, 8),
    to_signed(4, 8),
    to_signed(4, 8),
    to_signed(3, 8),
    to_signed(3, 8),
    to_signed(2, 8),
    to_signed(2, 8),
    to_signed(3, 8),
    to_signed(2, 8),
    to_signed(2, 8),
    to_signed(2, 8),
    to_signed(2, 8),
    to_signed(3, 8),
    to_signed(4, 8),
    to_signed(5, 8),
    to_signed(6, 8),
    to_signed(6, 8),
    to_signed(6, 8),
    to_signed(6, 8),
    to_signed(6, 8),
    to_signed(6, 8),
    to_signed(5, 8),
    to_signed(6, 8),
    to_signed(6, 8),
    to_signed(6, 8),
    to_signed(5, 8),
    to_signed(4, 8),
    to_signed(3, 8),
    to_signed(3, 8),
    to_signed(3, 8),
    to_signed(2, 8),
    to_signed(2, 8),
    to_signed(3, 8),
    to_signed(3, 8),
    to_signed(4, 8),
    to_signed(5, 8),
    to_signed(5, 8),
    to_signed(6, 8),
    to_signed(7, 8),
    to_signed(7, 8),
    to_signed(8, 8),
    to_signed(8, 8),
    to_signed(8, 8),
    to_signed(8, 8),
    to_signed(8, 8),
    to_signed(8, 8),
    to_signed(8, 8),
    to_signed(8, 8),
    to_signed(7, 8),
    to_signed(6, 8),
    to_signed(6, 8),
    to_signed(7, 8),
    to_signed(6, 8),
    to_signed(6, 8),
    to_signed(6, 8),
    to_signed(7, 8),
    to_signed(7, 8),
    to_signed(8, 8),
    to_signed(8, 8),
    to_signed(8, 8),
    to_signed(8, 8),
    to_signed(8, 8),
    to_signed(8, 8),
    to_signed(8, 8),
    to_signed(8, 8),
    to_signed(7, 8),
    to_signed(7, 8),
    to_signed(7, 8),
    to_signed(6, 8),
    to_signed(6, 8),
    to_signed(5, 8),
    to_signed(4, 8),
    to_signed(4, 8),
    to_signed(3, 8),
    to_signed(3, 8),
    to_signed(3, 8),
    to_signed(3, 8),
    to_signed(3, 8),
    to_signed(3, 8),
    to_signed(3, 8),
    to_signed(3, 8),
    to_signed(4, 8),
    to_signed(4, 8),
    to_signed(4, 8),
    to_signed(3, 8),
    to_signed(3, 8),
    to_signed(3, 8),
    to_signed(2, 8),
    to_signed(2, 8),
    to_signed(1, 8),
    to_signed(1, 8),
    to_signed(1, 8),
    to_signed(0, 8),
    to_signed(0, 8),
    to_signed(-1, 8),
    to_signed(-2, 8),
    to_signed(-2, 8),
    to_signed(-1, 8),
    to_signed(-1, 8),
    to_signed(-1, 8),
    to_signed(-1, 8),
    to_signed(-1, 8),
    to_signed(-1, 8),
    to_signed(0, 8),
    to_signed(1, 8),
    to_signed(0, 8),
    to_signed(0, 8),
    to_signed(0, 8),
    to_signed(-1, 8),
    to_signed(-2, 8),
    to_signed(-2, 8),
    to_signed(-3, 8),
    to_signed(-4, 8),
    to_signed(-4, 8),
    to_signed(-5, 8),
    to_signed(-6, 8),
    to_signed(-7, 8),
    to_signed(-7, 8),
    to_signed(-6, 8),
    to_signed(-6, 8),
    to_signed(-6, 8),
    to_signed(-6, 8),
    to_signed(-7, 8),
    to_signed(-7, 8),
    to_signed(-6, 8),
    to_signed(-5, 8),
    to_signed(-5, 8),
    to_signed(-5, 8),
    to_signed(-5, 8),
    to_signed(-5, 8),
    to_signed(-6, 8),
    to_signed(-7, 8),
    to_signed(-7, 8),
    to_signed(-7, 8),
    to_signed(-7, 8),
    to_signed(-8, 8),
    to_signed(-8, 8),
    to_signed(-9, 8),
    to_signed(-10, 8),
    to_signed(-11, 8),
    to_signed(-11, 8),
    to_signed(-11, 8),
    to_signed(-10, 8),
    to_signed(-10, 8),
    to_signed(-10, 8),
    to_signed(-10, 8),
    to_signed(-10, 8),
    to_signed(-9, 8),
    to_signed(-9, 8),
    to_signed(-9, 8),
    to_signed(-9, 8),
    to_signed(-10, 8),
    to_signed(-10, 8),
    to_signed(-11, 8),
    to_signed(-11, 8),
    to_signed(-12, 8),
    to_signed(-12, 8),
    to_signed(-13, 8),
    to_signed(-14, 8),
    to_signed(-15, 8),
    to_signed(-16, 8),
    to_signed(-16, 8),
    to_signed(-15, 8),
    to_signed(-14, 8),
    to_signed(-14, 8),
    to_signed(-13, 8),
    to_signed(-13, 8),
    to_signed(-13, 8),
    to_signed(-13, 8),
    to_signed(-12, 8),
    to_signed(-11, 8),
    to_signed(-10, 8),
    to_signed(-11, 8),
    to_signed(-11, 8),
    to_signed(-11, 8),
    to_signed(-11, 8),
    to_signed(-11, 8),
    to_signed(-11, 8),
    to_signed(-11, 8),
    to_signed(-11, 8),
    to_signed(-12, 8),
    to_signed(-13, 8),
    to_signed(-13, 8),
    to_signed(-13, 8),
    to_signed(-12, 8),
    to_signed(-11, 8),
    to_signed(-11, 8),
    to_signed(-10, 8),
    to_signed(-10, 8),
    to_signed(-10, 8),
    to_signed(-10, 8),
    to_signed(-9, 8),
    to_signed(-9, 8),
    to_signed(-8, 8),
    to_signed(-9, 8),
    to_signed(-9, 8),
    to_signed(-9, 8),
    to_signed(-9, 8),
    to_signed(-10, 8),
    to_signed(-11, 8),
    to_signed(-11, 8),
    to_signed(-11, 8),
    to_signed(-11, 8),
    to_signed(-12, 8),
    to_signed(-13, 8),
    to_signed(-13, 8),
    to_signed(-13, 8),
    to_signed(-12, 8),
    to_signed(-11, 8),
    to_signed(-11, 8),
    to_signed(-10, 8),
    to_signed(-10, 8),
    to_signed(-10, 8),
    to_signed(-8, 8),
    to_signed(-7, 8),
    to_signed(-6, 8),
    to_signed(-5, 8),
    to_signed(-5, 8),
    to_signed(-5, 8),
    to_signed(-5, 8),
    to_signed(-6, 8),
    to_signed(-6, 8),
    to_signed(-5, 8),
    to_signed(-5, 8),
    to_signed(-5, 8),
    to_signed(-5, 8),
    to_signed(-6, 8),
    to_signed(-6, 8),
    to_signed(-5, 8),
    to_signed(-3, 8),
    to_signed(-2, 8),
    to_signed(-2, 8),
    to_signed(-1, 8),
    to_signed(-1, 8),
    to_signed(0, 8),
    to_signed(0, 8),
    to_signed(1, 8),
    to_signed(2, 8),
    to_signed(2, 8),
    to_signed(2, 8),
    to_signed(2, 8),
    to_signed(1, 8),
    to_signed(1, 8),
    to_signed(1, 8),
    to_signed(0, 8),
    to_signed(0, 8),
    to_signed(-1, 8),
    to_signed(-2, 8),
    to_signed(-3, 8),
    to_signed(-3, 8),
    to_signed(-2, 8),
    to_signed(0, 8),
    to_signed(0, 8),
    to_signed(0, 8),
    to_signed(0, 8),
    to_signed(0, 8),
    to_signed(0, 8),
    to_signed(1, 8),
    to_signed(2, 8),
    to_signed(2, 8),
    to_signed(3, 8),
    to_signed(2, 8),
    to_signed(2, 8),
    to_signed(1, 8),
    to_signed(1, 8),
    to_signed(1, 8),
    to_signed(1, 8),
    to_signed(1, 8),
    to_signed(1, 8),
    to_signed(0, 8),
    to_signed(0, 8),
    to_signed(0, 8),
    to_signed(2, 8),
    to_signed(3, 8),
    to_signed(5, 8),
    to_signed(5, 8),
    to_signed(6, 8),
    to_signed(6, 8),
    to_signed(7, 8),
    to_signed(8, 8),
    to_signed(9, 8),
    to_signed(10, 8),
    to_signed(10, 8),
    to_signed(10, 8),
    to_signed(9, 8),
    to_signed(9, 8),
    to_signed(8, 8),
    to_signed(7, 8),
    to_signed(7, 8),
    to_signed(7, 8),
    to_signed(6, 8),
    to_signed(6, 8),
    to_signed(5, 8),
    to_signed(4, 8),
    to_signed(5, 8),
    to_signed(5, 8),
    to_signed(5, 8),
    to_signed(5, 8),
    to_signed(5, 8),
    to_signed(4, 8),
    to_signed(4, 8),
    to_signed(5, 8),
    to_signed(5, 8),
    to_signed(5, 8),
    to_signed(5, 8),
    to_signed(4, 8),
    to_signed(3, 8),
    to_signed(2, 8),
    to_signed(1, 8),
    to_signed(1, 8),
    to_signed(0, 8),
    to_signed(0, 8),
    to_signed(-1, 8),
    to_signed(-2, 8),
    to_signed(-3, 8),
    to_signed(-3, 8),
    to_signed(-2, 8),
    to_signed(-1, 8),
    to_signed(0, 8),
    to_signed(0, 8),
    to_signed(0, 8),
    to_signed(0, 8),
    to_signed(0, 8),
    to_signed(1, 8),
    to_signed(1, 8),
    to_signed(2, 8),
    to_signed(2, 8),
    to_signed(3, 8),
    to_signed(3, 8),
    to_signed(3, 8),
    to_signed(3, 8),
    to_signed(2, 8),
    to_signed(3, 8),
    to_signed(3, 8),
    to_signed(3, 8),
    to_signed(2, 8),
    to_signed(1, 8),
    to_signed(1, 8),
    to_signed(2, 8),
    to_signed(4, 8),
    to_signed(5, 8),
    to_signed(5, 8),
    to_signed(4, 8),
    to_signed(4, 8),
    to_signed(4, 8),
    to_signed(5, 8),
    to_signed(5, 8),
    to_signed(6, 8),
    to_signed(6, 8),
    to_signed(6, 8),
    to_signed(7, 8),
    to_signed(6, 8),
    to_signed(6, 8),
    to_signed(5, 8),
    to_signed(5, 8),
    to_signed(5, 8),
    to_signed(5, 8),
    to_signed(4, 8),
    to_signed(3, 8),
    to_signed(3, 8),
    to_signed(3, 8),
    to_signed(4, 8),
    to_signed(5, 8),
    to_signed(5, 8),
    to_signed(5, 8),
    to_signed(4, 8),
    to_signed(4, 8),
    to_signed(4, 8),
    to_signed(4, 8),
    to_signed(4, 8),
    to_signed(4, 8),
    to_signed(4, 8),
    to_signed(4, 8),
    to_signed(3, 8),
    to_signed(2, 8),
    to_signed(1, 8),
    to_signed(0, 8),
    to_signed(0, 8),
    to_signed(-1, 8),
    to_signed(-2, 8),
    to_signed(-2, 8),
    to_signed(-2, 8),
    to_signed(-1, 8),
    to_signed(-1, 8),
    to_signed(0, 8),
    to_signed(0, 8),
    to_signed(1, 8),
    to_signed(1, 8),
    to_signed(1, 8),
    to_signed(1, 8),
    to_signed(1, 8),
    to_signed(2, 8),
    to_signed(3, 8),
    to_signed(3, 8),
    to_signed(3, 8),
    to_signed(3, 8),
    to_signed(2, 8),
    to_signed(1, 8),
    to_signed(0, 8),
    to_signed(1, 8),
    to_signed(1, 8),
    to_signed(1, 8),
    to_signed(0, 8),
    to_signed(0, 8),
    to_signed(1, 8),
    to_signed(3, 8),
    to_signed(4, 8),
    to_signed(4, 8),
    to_signed(3, 8),
    to_signed(3, 8),
    to_signed(3, 8),
    to_signed(3, 8),
    to_signed(2, 8),
    to_signed(1, 8),
    to_signed(1, 8),
    to_signed(0, 8),
    to_signed(0, 8),
    to_signed(0, 8),
    to_signed(-1, 8),
    to_signed(-3, 8),
    to_signed(-4, 8),
    to_signed(-4, 8),
    to_signed(-5, 8),
    to_signed(-6, 8),
    to_signed(-7, 8),
    to_signed(-7, 8),
    to_signed(-7, 8),
    to_signed(-6, 8),
    to_signed(-5, 8),
    to_signed(-5, 8),
    to_signed(-5, 8),
    to_signed(-5, 8),
    to_signed(-4, 8),
    to_signed(-4, 8),
    to_signed(-4, 8),
    to_signed(-4, 8),
    to_signed(-4, 8),
    to_signed(-4, 8),
    to_signed(-4, 8),
    to_signed(-4, 8),
    to_signed(-4, 8),
    to_signed(-4, 8),
    to_signed(-5, 8),
    to_signed(-5, 8),
    to_signed(-6, 8),
    to_signed(-6, 8),
    to_signed(-6, 8),
    to_signed(-5, 8),
    to_signed(-4, 8),
    to_signed(-3, 8),
    to_signed(-2, 8),
    to_signed(-2, 8),
    to_signed(-2, 8),
    to_signed(-2, 8),
    to_signed(-1, 8),
    to_signed(-1, 8),
    to_signed(-1, 8),
    to_signed(-1, 8),
    to_signed(-1, 8),
    to_signed(-1, 8),
    to_signed(0, 8),
    to_signed(0, 8),
    to_signed(-1, 8),
    to_signed(-2, 8),
    to_signed(-3, 8),
    to_signed(-4, 8),
    to_signed(-4, 8),
    to_signed(-5, 8),
    to_signed(-5, 8),
    to_signed(-5, 8),
    to_signed(-4, 8),
    to_signed(-3, 8),
    to_signed(-2, 8),
    to_signed(-1, 8),
    to_signed(-1, 8),
    to_signed(0, 8),
    to_signed(0, 8),
    to_signed(1, 8),
    to_signed(1, 8),
    to_signed(0, 8),
    to_signed(1, 8),
    to_signed(1, 8),
    to_signed(1, 8),
    to_signed(1, 8),
    to_signed(1, 8),
    to_signed(0, 8),
    to_signed(0, 8),
    to_signed(0, 8),
    to_signed(0, 8),
    to_signed(0, 8),
    to_signed(0, 8),
    to_signed(0, 8),
    to_signed(1, 8),
    to_signed(2, 8),
    to_signed(3, 8),
    to_signed(4, 8),
    to_signed(4, 8),
    to_signed(4, 8),
    to_signed(5, 8),
    to_signed(5, 8),
    to_signed(5, 8),
    to_signed(4, 8),
    to_signed(4, 8),
    to_signed(4, 8),
    to_signed(5, 8),
    to_signed(5, 8),
    to_signed(4, 8),
    to_signed(4, 8),
    to_signed(3, 8),
    to_signed(2, 8),
    to_signed(2, 8),
    to_signed(2, 8),
    to_signed(2, 8),
    to_signed(2, 8),
    to_signed(2, 8),
    to_signed(2, 8),
    to_signed(3, 8),
    to_signed(4, 8),
    to_signed(4, 8),
    to_signed(4, 8),
    to_signed(4, 8),
    to_signed(4, 8),
    to_signed(4, 8),
    to_signed(4, 8),
    to_signed(4, 8),
    to_signed(4, 8),
    to_signed(5, 8),
    to_signed(5, 8),
    to_signed(4, 8),
    to_signed(4, 8),
    to_signed(3, 8),
    to_signed(3, 8),
    to_signed(3, 8),
    to_signed(3, 8),
    to_signed(3, 8),
    to_signed(3, 8),
    to_signed(4, 8),
    to_signed(5, 8),
    to_signed(5, 8),
    to_signed(5, 8),
    to_signed(5, 8),
    to_signed(5, 8),
    to_signed(6, 8),
    to_signed(6, 8),
    to_signed(6, 8),
    to_signed(5, 8),
    to_signed(5, 8),
    to_signed(5, 8),
    to_signed(5, 8),
    to_signed(4, 8),
    to_signed(4, 8),
    to_signed(3, 8),
    to_signed(2, 8),
    to_signed(1, 8),
    to_signed(1, 8),
    to_signed(0, 8),
    to_signed(-1, 8),
    to_signed(-1, 8),
    to_signed(0, 8),
    to_signed(1, 8),
    to_signed(1, 8),
    to_signed(0, 8),
    to_signed(0, 8),
    to_signed(0, 8),
    to_signed(0, 8),
    to_signed(1, 8),
    to_signed(0, 8),
    to_signed(0, 8),
    to_signed(-1, 8),
    to_signed(-1, 8),
    to_signed(-1, 8),
    to_signed(-1, 8),
    to_signed(-1, 8),
    to_signed(-2, 8),
    to_signed(-2, 8),
    to_signed(-3, 8),
    to_signed(-4, 8),
    to_signed(-4, 8),
    to_signed(-4, 8),
    to_signed(-4, 8),
    to_signed(-3, 8),
    to_signed(-1, 8),
    to_signed(-1, 8),
    to_signed(0, 8),
    to_signed(0, 8),
    to_signed(0, 8),
    to_signed(1, 8),
    to_signed(2, 8),
    to_signed(1, 8),
    to_signed(1, 8),
    to_signed(1, 8),
    to_signed(1, 8),
    to_signed(2, 8),
    to_signed(2, 8),
    to_signed(1, 8),
    to_signed(1, 8),
    to_signed(1, 8),
    to_signed(1, 8),
    to_signed(0, 8),
    to_signed(-1, 8),
    to_signed(-1, 8),
    to_signed(0, 8),
    to_signed(1, 8),
    to_signed(2, 8),
    to_signed(2, 8),
    to_signed(2, 8),
    to_signed(2, 8),
    to_signed(2, 8),
    to_signed(3, 8),
    to_signed(3, 8),
    to_signed(2, 8),
    to_signed(2, 8),
    to_signed(2, 8),
    to_signed(1, 8),
    to_signed(1, 8),
    to_signed(0, 8),
    to_signed(0, 8),
    to_signed(0, 8),
    to_signed(0, 8),
    to_signed(-1, 8),
    to_signed(-2, 8),
    to_signed(-3, 8),
    to_signed(-3, 8),
    to_signed(-3, 8),
    to_signed(-2, 8),
    to_signed(-2, 8),
    to_signed(-1, 8),
    to_signed(-1, 8),
    to_signed(0, 8),
    to_signed(0, 8),
    to_signed(1, 8),
    to_signed(1, 8),
    to_signed(1, 8),
    to_signed(0, 8),
    to_signed(0, 8),
    to_signed(0, 8),
    to_signed(0, 8),
    to_signed(0, 8),
    to_signed(0, 8),
    to_signed(1, 8),
    to_signed(1, 8),
    to_signed(1, 8),
    to_signed(0, 8),
    to_signed(0, 8),
    to_signed(0, 8),
    to_signed(0, 8),
    to_signed(1, 8),
    to_signed(2, 8),
    to_signed(2, 8),
    to_signed(3, 8),
    to_signed(3, 8),
    to_signed(3, 8),
    to_signed(4, 8),
    to_signed(4, 8),
    to_signed(4, 8),
    to_signed(3, 8),
    to_signed(3, 8),
    to_signed(2, 8),
    to_signed(2, 8),
    to_signed(2, 8),
    to_signed(2, 8),
    to_signed(2, 8),
    to_signed(1, 8),
    to_signed(0, 8),
    to_signed(0, 8),
    to_signed(-1, 8),
    to_signed(-2, 8),
    to_signed(-2, 8),
    to_signed(-2, 8),
    to_signed(-1, 8),
    to_signed(-1, 8),
    to_signed(-1, 8),
    to_signed(0, 8),
    to_signed(0, 8),
    to_signed(0, 8),
    to_signed(1, 8),
    to_signed(0, 8),
    to_signed(0, 8),
    to_signed(0, 8),
    to_signed(0, 8),
    to_signed(0, 8),
    to_signed(0, 8),
    to_signed(0, 8),
    to_signed(0, 8),
    to_signed(0, 8),
    to_signed(-1, 8),
    to_signed(-1, 8),
    to_signed(-1, 8),
    to_signed(-2, 8),
    to_signed(-2, 8),
    to_signed(-1, 8),
    to_signed(0, 8),
    to_signed(1, 8),
    to_signed(1, 8),
    to_signed(1, 8),
    to_signed(1, 8),
    to_signed(1, 8),
    to_signed(2, 8),
    to_signed(1, 8),
    to_signed(1, 8),
    to_signed(0, 8),
    to_signed(0, 8),
    to_signed(-1, 8),
    to_signed(-1, 8),
    to_signed(-2, 8),
    to_signed(-2, 8),
    to_signed(-3, 8),
    to_signed(-3, 8),
    to_signed(-4, 8),
    to_signed(-5, 8),
    to_signed(-6, 8),
    to_signed(-7, 8),
    to_signed(-6, 8),
    to_signed(-5, 8),
    to_signed(-4, 8),
    to_signed(-4, 8),
    to_signed(-5, 8),
    to_signed(-5, 8),
    to_signed(-4, 8),
    to_signed(-4, 8),
    to_signed(-4, 8),
    to_signed(-4, 8),
    to_signed(-5, 8),
    to_signed(-5, 8),
    to_signed(-6, 8),
    to_signed(-6, 8),
    to_signed(-6, 8),
    to_signed(-6, 8),
    to_signed(-6, 8),
    to_signed(-5, 8),
    to_signed(-5, 8),
    to_signed(-5, 8),
    to_signed(-6, 8),
    to_signed(-6, 8),
    to_signed(-4, 8),
    to_signed(-3, 8),
    to_signed(-2, 8),
    to_signed(-1, 8),
    to_signed(-1, 8),
    to_signed(-1, 8),
    to_signed(0, 8),
    to_signed(0, 8),
    to_signed(1, 8),
    to_signed(1, 8),
    to_signed(1, 8),
    to_signed(1, 8),
    to_signed(0, 8),
    to_signed(-1, 8),
    to_signed(-1, 8),
    to_signed(-1, 8),
    to_signed(-1, 8),
    to_signed(-1, 8),
    to_signed(-1, 8),
    to_signed(-2, 8),
    to_signed(-3, 8),
    to_signed(-3, 8),
    to_signed(-3, 8),
    to_signed(-2, 8),
    to_signed(-1, 8),
    to_signed(-1, 8),
    to_signed(-2, 8),
    to_signed(-2, 8),
    to_signed(-2, 8),
    to_signed(-3, 8),
    to_signed(-3, 8),
    to_signed(-3, 8),
    to_signed(-3, 8),
    to_signed(-4, 8),
    to_signed(-5, 8),
    to_signed(-6, 8),
    to_signed(-6, 8),
    to_signed(-6, 8),
    to_signed(-5, 8),
    to_signed(-5, 8),
    to_signed(-6, 8),
    to_signed(-6, 8),
    to_signed(-6, 8),
    to_signed(-7, 8),
    to_signed(-6, 8),
    to_signed(-5, 8),
    to_signed(-4, 8),
    to_signed(-3, 8),
    to_signed(-3, 8),
    to_signed(-3, 8),
    to_signed(-3, 8),
    to_signed(-2, 8),
    to_signed(-2, 8),
    to_signed(-1, 8),
    to_signed(0, 8),
    to_signed(0, 8),
    to_signed(-1, 8),
    to_signed(-1, 8),
    to_signed(-1, 8),
    to_signed(-1, 8),
    to_signed(0, 8),
    to_signed(0, 8),
    to_signed(-1, 8),
    to_signed(-2, 8),
    to_signed(-2, 8),
    to_signed(-2, 8),
    to_signed(-2, 8),
    to_signed(-1, 8),
    to_signed(0, 8),
    to_signed(1, 8),
    to_signed(1, 8),
    to_signed(0, 8),
    to_signed(-1, 8),
    to_signed(-1, 8),
    to_signed(0, 8),
    to_signed(0, 8),
    to_signed(0, 8),
    to_signed(-1, 8),
    to_signed(-2, 8),
    to_signed(-2, 8),
    to_signed(-3, 8),
    to_signed(-2, 8),
    to_signed(-2, 8),
    to_signed(-2, 8),
    to_signed(-3, 8),
    to_signed(-4, 8),
    to_signed(-5, 8),
    to_signed(-5, 8),
    to_signed(-4, 8),
    to_signed(-3, 8),
    to_signed(-2, 8),
    to_signed(-2, 8),
    to_signed(-1, 8),
    to_signed(-1, 8),
    to_signed(-2, 8),
    to_signed(-2, 8),
    to_signed(-1, 8),
    to_signed(0, 8),
    to_signed(1, 8),
    to_signed(1, 8),
    to_signed(0, 8),
    to_signed(0, 8),
    to_signed(0, 8),
    to_signed(1, 8),
    to_signed(1, 8),
    to_signed(1, 8),
    to_signed(0, 8),
    to_signed(0, 8),
    to_signed(-1, 8),
    to_signed(-1, 8),
    to_signed(0, 8),
    to_signed(0, 8),
    to_signed(2, 8),
    to_signed(3, 8),
    to_signed(3, 8),
    to_signed(3, 8),
    to_signed(2, 8),
    to_signed(2, 8),
    to_signed(3, 8),
    to_signed(3, 8),
    to_signed(3, 8),
    to_signed(3, 8),
    to_signed(2, 8),
    to_signed(1, 8),
    to_signed(0, 8),
    to_signed(0, 8),
    to_signed(1, 8),
    to_signed(2, 8),
    to_signed(0, 8),
    to_signed(-2, 8),
    to_signed(-3, 8),
    to_signed(-2, 8),
    to_signed(-1, 8),
    to_signed(0, 8),
    to_signed(1, 8),
    to_signed(1, 8),
    to_signed(1, 8),
    to_signed(1, 8),
    to_signed(1, 8),
    to_signed(2, 8),
    to_signed(3, 8),
    to_signed(3, 8),
    to_signed(4, 8),
    to_signed(4, 8),
    to_signed(4, 8),
    to_signed(4, 8),
    to_signed(3, 8),
    to_signed(4, 8),
    to_signed(4, 8),
    to_signed(5, 8),
    to_signed(4, 8),
    to_signed(3, 8),
    to_signed(2, 8),
    to_signed(2, 8),
    to_signed(3, 8),
    to_signed(5, 8),
    to_signed(6, 8),
    to_signed(7, 8),
    to_signed(6, 8),
    to_signed(6, 8),
    to_signed(6, 8),
    to_signed(6, 8),
    to_signed(6, 8),
    to_signed(7, 8),
    to_signed(7, 8),
    to_signed(6, 8),
    to_signed(5, 8),
    to_signed(4, 8),
    to_signed(3, 8),
    to_signed(4, 8),
    to_signed(3, 8),
    to_signed(3, 8),
    to_signed(2, 8),
    to_signed(0, 8),
    to_signed(-1, 8),
    to_signed(-1, 8),
    to_signed(-1, 8),
    to_signed(0, 8),
    to_signed(1, 8),
    to_signed(1, 8),
    to_signed(1, 8),
    to_signed(1, 8),
    to_signed(1, 8),
    to_signed(0, 8),
    to_signed(1, 8),
    to_signed(1, 8),
    to_signed(1, 8),
    to_signed(1, 8),
    to_signed(1, 8),
    to_signed(0, 8),
    to_signed(0, 8),
    to_signed(0, 8),
    to_signed(1, 8),
    to_signed(1, 8),
    to_signed(1, 8),
    to_signed(1, 8),
    to_signed(0, 8),
    to_signed(0, 8),
    to_signed(1, 8),
    to_signed(2, 8),
    to_signed(3, 8),
    to_signed(4, 8),
    to_signed(4, 8),
    to_signed(4, 8),
    to_signed(4, 8),
    to_signed(4, 8),
    to_signed(4, 8),
    to_signed(6, 8),
    to_signed(6, 8),
    to_signed(6, 8),
    to_signed(5, 8),
    to_signed(5, 8),
    to_signed(4, 8),
    to_signed(4, 8),
    to_signed(5, 8),
    to_signed(4, 8),
    to_signed(4, 8),
    to_signed(3, 8),
    to_signed(2, 8),
    to_signed(1, 8),
    to_signed(1, 8),
    to_signed(2, 8),
    to_signed(3, 8),
    to_signed(4, 8),
    to_signed(4, 8),
    to_signed(3, 8),
    to_signed(1, 8),
    to_signed(1, 8),
    to_signed(1, 8),
    to_signed(1, 8),
    to_signed(1, 8),
    to_signed(1, 8),
    to_signed(0, 8),
    to_signed(-1, 8),
    to_signed(-2, 8),
    to_signed(-2, 8),
    to_signed(-2, 8),
    to_signed(-2, 8),
    to_signed(-3, 8),
    to_signed(-4, 8),
    to_signed(-5, 8),
    to_signed(-5, 8),
    to_signed(-5, 8),
    to_signed(-4, 8),
    to_signed(-3, 8),
    to_signed(-2, 8),
    to_signed(-2, 8),
    to_signed(-3, 8),
    to_signed(-3, 8),
    to_signed(-3, 8),
    to_signed(-2, 8),
    to_signed(-1, 8),
    to_signed(-1, 8),
    to_signed(-1, 8),
    to_signed(-1, 8),
    to_signed(-2, 8),
    to_signed(-2, 8),
    to_signed(-1, 8),
    to_signed(0, 8),
    to_signed(0, 8),
    to_signed(-1, 8),
    to_signed(-1, 8),
    to_signed(-2, 8),
    to_signed(-2, 8),
    to_signed(-1, 8),
    to_signed(0, 8),
    to_signed(0, 8),
    to_signed(1, 8),
    to_signed(1, 8),
    to_signed(1, 8),
    to_signed(0, 8),
    to_signed(0, 8),
    to_signed(0, 8),
    to_signed(1, 8),
    to_signed(1, 8),
    to_signed(1, 8),
    to_signed(1, 8),
    to_signed(0, 8),
    to_signed(-1, 8),
    to_signed(-1, 8),
    to_signed(0, 8),
    to_signed(0, 8),
    to_signed(-1, 8),
    to_signed(-2, 8),
    to_signed(-3, 8),
    to_signed(-3, 8),
    to_signed(-3, 8),
    to_signed(-2, 8),
    to_signed(-1, 8),
    to_signed(-1, 8),
    to_signed(-1, 8),
    to_signed(-1, 8),
    to_signed(-2, 8),
    to_signed(-2, 8),
    to_signed(-1, 8),
    to_signed(-1, 8),
    to_signed(0, 8),
    to_signed(-1, 8),
    to_signed(-1, 8),
    to_signed(-1, 8),
    to_signed(-1, 8),
    to_signed(-2, 8),
    to_signed(-2, 8),
    to_signed(-2, 8),
    to_signed(-1, 8),
    to_signed(-1, 8),
    to_signed(-2, 8),
    to_signed(-2, 8),
    to_signed(-2, 8),
    to_signed(-1, 8),
    to_signed(0, 8),
    to_signed(1, 8),
    to_signed(1, 8),
    to_signed(1, 8),
    to_signed(0, 8),
    to_signed(0, 8),
    to_signed(1, 8),
    to_signed(1, 8),
    to_signed(2, 8),
    to_signed(2, 8),
    to_signed(1, 8),
    to_signed(0, 8),
    to_signed(0, 8),
    to_signed(0, 8),
    to_signed(0, 8),
    to_signed(0, 8),
    to_signed(-1, 8),
    to_signed(-2, 8),
    to_signed(-3, 8),
    to_signed(-4, 8),
    to_signed(-4, 8),
    to_signed(-3, 8),
    to_signed(-3, 8),
    to_signed(-2, 8),
    to_signed(-2, 8),
    to_signed(-3, 8),
    to_signed(-3, 8),
    to_signed(-3, 8),
    to_signed(-3, 8),
    to_signed(-3, 8),
    to_signed(-3, 8),
    to_signed(-3, 8),
    to_signed(-4, 8),
    to_signed(-4, 8),
    to_signed(-5, 8),
    to_signed(-5, 8),
    to_signed(-5, 8),
    to_signed(-5, 8),
    to_signed(-5, 8),
    to_signed(-6, 8),
    to_signed(-7, 8),
    to_signed(-7, 8),
    to_signed(-8, 8),
    to_signed(-7, 8),
    to_signed(-6, 8),
    to_signed(-5, 8),
    to_signed(-5, 8),
    to_signed(-5, 8),
    to_signed(-5, 8),
    to_signed(-4, 8),
    to_signed(-4, 8),
    to_signed(-3, 8),
    to_signed(-3, 8),
    to_signed(-3, 8),
    to_signed(-3, 8),
    to_signed(-3, 8),
    to_signed(-4, 8),
    to_signed(-4, 8),
    to_signed(-3, 8),
    to_signed(-3, 8),
    to_signed(-4, 8),
    to_signed(-5, 8),
    to_signed(-5, 8),
    to_signed(-5, 8),
    to_signed(-5, 8),
    to_signed(-5, 8),
    to_signed(-4, 8),
    to_signed(-4, 8),
    to_signed(-4, 8),
    to_signed(-4, 8),
    to_signed(-4, 8),
    to_signed(-4, 8),
    to_signed(-4, 8),
    to_signed(-4, 8),
    to_signed(-4, 8),
    to_signed(-4, 8),
    to_signed(-4, 8),
    to_signed(-4, 8),
    to_signed(-4, 8),
    to_signed(-4, 8),
    to_signed(-4, 8),
    to_signed(-4, 8),
    to_signed(-4, 8),
    to_signed(-3, 8),
    to_signed(-3, 8),
    to_signed(-4, 8),
    to_signed(-3, 8),
    to_signed(-3, 8),
    to_signed(-2, 8),
    to_signed(-1, 8),
    to_signed(-1, 8),
    to_signed(-1, 8),
    to_signed(-1, 8),
    to_signed(0, 8),
    to_signed(0, 8),
    to_signed(1, 8),
    to_signed(1, 8),
    to_signed(1, 8),
    to_signed(1, 8),
    to_signed(1, 8),
    to_signed(1, 8),
    to_signed(0, 8),
    to_signed(0, 8),
    to_signed(0, 8),
    to_signed(0, 8),
    to_signed(-1, 8),
    to_signed(-1, 8),
    to_signed(-2, 8),
    to_signed(-2, 8),
    to_signed(-2, 8),
    to_signed(-1, 8),
    to_signed(-2, 8),
    to_signed(-2, 8),
    to_signed(-3, 8),
    to_signed(-3, 8),
    to_signed(-3, 8),
    to_signed(-3, 8),
    to_signed(-3, 8),
    to_signed(-4, 8),
    to_signed(-4, 8),
    to_signed(-4, 8),
    to_signed(-4, 8),
    to_signed(-5, 8),
    to_signed(-6, 8),
    to_signed(-6, 8),
    to_signed(-5, 8),
    to_signed(-5, 8),
    to_signed(-5, 8),
    to_signed(-6, 8),
    to_signed(-6, 8),
    to_signed(-5, 8),
    to_signed(-5, 8),
    to_signed(-4, 8),
    to_signed(-3, 8),
    to_signed(-3, 8),
    to_signed(-2, 8),
    to_signed(-2, 8),
    to_signed(-2, 8),
    to_signed(-1, 8),
    to_signed(-1, 8),
    to_signed(-1, 8),
    to_signed(0, 8),
    to_signed(0, 8),
    to_signed(0, 8),
    to_signed(0, 8),
    to_signed(0, 8),
    to_signed(0, 8),
    to_signed(1, 8),
    to_signed(1, 8),
    to_signed(1, 8),
    to_signed(1, 8),
    to_signed(1, 8),
    to_signed(1, 8),
    to_signed(1, 8),
    to_signed(1, 8),
    to_signed(2, 8),
    to_signed(2, 8),
    to_signed(2, 8),
    to_signed(2, 8),
    to_signed(2, 8),
    to_signed(2, 8),
    to_signed(2, 8),
    to_signed(2, 8),
    to_signed(2, 8),
    to_signed(2, 8),
    to_signed(2, 8),
    to_signed(1, 8),
    to_signed(0, 8),
    to_signed(-1, 8),
    to_signed(-1, 8),
    to_signed(0, 8),
    to_signed(0, 8),
    to_signed(-1, 8),
    to_signed(-1, 8),
    to_signed(-1, 8),
    to_signed(-1, 8),
    to_signed(-1, 8),
    to_signed(0, 8),
    to_signed(-1, 8),
    to_signed(0, 8),
    to_signed(0, 8),
    to_signed(1, 8),
    to_signed(2, 8),
    to_signed(2, 8),
    to_signed(2, 8),
    to_signed(2, 8),
    to_signed(2, 8),
    to_signed(2, 8),
    to_signed(2, 8),
    to_signed(1, 8),
    to_signed(1, 8),
    to_signed(1, 8),
    to_signed(2, 8),
    to_signed(2, 8),
    to_signed(2, 8),
    to_signed(1, 8),
    to_signed(1, 8),
    to_signed(1, 8),
    to_signed(2, 8),
    to_signed(2, 8),
    to_signed(2, 8),
    to_signed(2, 8),
    to_signed(3, 8),
    to_signed(4, 8),
    to_signed(4, 8),
    to_signed(4, 8),
    to_signed(4, 8),
    to_signed(5, 8),
    to_signed(5, 8),
    to_signed(5, 8),
    to_signed(4, 8),
    to_signed(4, 8),
    to_signed(3, 8),
    to_signed(4, 8),
    to_signed(4, 8),
    to_signed(4, 8),
    to_signed(3, 8),
    to_signed(3, 8),
    to_signed(3, 8),
    to_signed(3, 8),
    to_signed(3, 8),
    to_signed(3, 8),
    to_signed(3, 8),
    to_signed(4, 8),
    to_signed(4, 8),
    to_signed(5, 8),
    to_signed(5, 8),
    to_signed(5, 8),
    to_signed(5, 8),
    to_signed(6, 8),
    to_signed(6, 8),
    to_signed(6, 8),
    to_signed(5, 8),
    to_signed(4, 8),
    to_signed(4, 8),
    to_signed(4, 8),
    to_signed(3, 8),
    to_signed(3, 8),
    to_signed(2, 8),
    to_signed(2, 8),
    to_signed(2, 8),
    to_signed(2, 8),
    to_signed(2, 8),
    to_signed(1, 8),
    to_signed(2, 8),
    to_signed(2, 8),
    to_signed(2, 8),
    to_signed(2, 8),
    to_signed(2, 8),
    to_signed(3, 8),
    to_signed(2, 8),
    to_signed(2, 8),
    to_signed(2, 8),
    to_signed(2, 8),
    to_signed(1, 8),
    to_signed(0, 8),
    to_signed(0, 8),
    to_signed(0, 8),
    to_signed(0, 8),
    to_signed(0, 8),
    to_signed(-1, 8),
    to_signed(-1, 8),
    to_signed(-1, 8),
    to_signed(-1, 8),
    to_signed(-1, 8),
    to_signed(-1, 8),
    to_signed(-2, 8),
    to_signed(-1, 8),
    to_signed(0, 8),
    to_signed(1, 8),
    to_signed(1, 8),
    to_signed(2, 8),
    to_signed(2, 8),
    to_signed(2, 8),
    to_signed(2, 8),
    to_signed(1, 8),
    to_signed(1, 8),
    to_signed(0, 8),
    to_signed(0, 8),
    to_signed(1, 8),
    to_signed(1, 8),
    to_signed(0, 8),
    to_signed(0, 8),
    to_signed(0, 8),
    to_signed(0, 8),
    to_signed(0, 8),
    to_signed(0, 8),
    to_signed(0, 8),
    to_signed(0, 8),
    to_signed(0, 8),
    to_signed(1, 8),
    to_signed(2, 8),
    to_signed(2, 8),
    to_signed(2, 8),
    to_signed(2, 8),
    to_signed(2, 8),
    to_signed(2, 8),
    to_signed(1, 8),
    to_signed(1, 8),
    to_signed(0, 8),
    to_signed(-1, 8),
    to_signed(0, 8),
    to_signed(0, 8),
    to_signed(0, 8),
    to_signed(0, 8),
    to_signed(-1, 8),
    to_signed(-1, 8),
    to_signed(-1, 8),
    to_signed(-2, 8),
    to_signed(-2, 8),
    to_signed(-2, 8),
    to_signed(-2, 8),
    to_signed(-1, 8),
    to_signed(-1, 8),
    to_signed(-1, 8),
    to_signed(-1, 8),
    to_signed(-1, 8),
    to_signed(0, 8),
    to_signed(0, 8),
    to_signed(-1, 8),
    to_signed(-2, 8),
    to_signed(-3, 8),
    to_signed(-3, 8),
    to_signed(-3, 8),
    to_signed(-2, 8),
    to_signed(-2, 8),
    to_signed(-2, 8),
    to_signed(-3, 8),
    to_signed(-3, 8),
    to_signed(-3, 8),
    to_signed(-3, 8),
    to_signed(-4, 8),
    to_signed(-4, 8),
    to_signed(-3, 8),
    to_signed(-3, 8),
    to_signed(-2, 8),
    to_signed(-2, 8),
    to_signed(-1, 8),
    to_signed(-1, 8),
    to_signed(0, 8),
    to_signed(-1, 8),
    to_signed(-1, 8),
    to_signed(-2, 8),
    to_signed(-3, 8),
    to_signed(-3, 8),
    to_signed(-2, 8),
    to_signed(-2, 8),
    to_signed(-2, 8),
    to_signed(-2, 8),
    to_signed(-2, 8),
    to_signed(-1, 8),
    to_signed(-2, 8),
    to_signed(-2, 8),
    to_signed(-3, 8),
    to_signed(-2, 8),
    to_signed(-1, 8),
    to_signed(0, 8),
    to_signed(1, 8),
    to_signed(1, 8),
    to_signed(1, 8),
    to_signed(2, 8),
    to_signed(2, 8),
    to_signed(3, 8),
    to_signed(2, 8),
    to_signed(2, 8),
    to_signed(2, 8),
    to_signed(3, 8),
    to_signed(4, 8),
    to_signed(4, 8),
    to_signed(4, 8),
    to_signed(4, 8),
    to_signed(5, 8),
    to_signed(5, 8),
    to_signed(5, 8),
    to_signed(4, 8),
    to_signed(3, 8),
    to_signed(4, 8),
    to_signed(4, 8),
    to_signed(5, 8),
    to_signed(5, 8),
    to_signed(5, 8),
    to_signed(6, 8),
    to_signed(6, 8),
    to_signed(6, 8),
    to_signed(5, 8),
    to_signed(5, 8),
    to_signed(3, 8),
    to_signed(2, 8),
    to_signed(2, 8),
    to_signed(1, 8),
    to_signed(1, 8),
    to_signed(0, 8),
    to_signed(0, 8),
    to_signed(0, 8),
    to_signed(-1, 8),
    to_signed(-1, 8),
    to_signed(-3, 8),
    to_signed(-3, 8),
    to_signed(-3, 8),
    to_signed(-3, 8),
    to_signed(-3, 8),
    to_signed(-3, 8),
    to_signed(-3, 8),
    to_signed(-2, 8),
    to_signed(-2, 8),
    to_signed(-1, 8),
    to_signed(-1, 8),
    to_signed(-2, 8),
    to_signed(-3, 8),
    to_signed(-3, 8),
    to_signed(-3, 8),
    to_signed(-2, 8),
    to_signed(-2, 8),
    to_signed(-2, 8),
    to_signed(-2, 8),
    to_signed(-1, 8),
    to_signed(-1, 8),
    to_signed(-1, 8),
    to_signed(-1, 8),
    to_signed(-2, 8),
    to_signed(-2, 8),
    to_signed(-1, 8),
    to_signed(0, 8),
    to_signed(1, 8),
    to_signed(1, 8),
    to_signed(2, 8),
    to_signed(2, 8),
    to_signed(3, 8),
    to_signed(3, 8),
    to_signed(3, 8),
    to_signed(2, 8),
    to_signed(1, 8),
    to_signed(1, 8),
    to_signed(1, 8),
    to_signed(1, 8),
    to_signed(1, 8),
    to_signed(0, 8),
    to_signed(0, 8),
    to_signed(0, 8),
    to_signed(-1, 8),
    to_signed(-2, 8),
    to_signed(-2, 8),
    to_signed(-2, 8),
    to_signed(-1, 8),
    to_signed(-1, 8),
    to_signed(-1, 8),
    to_signed(-1, 8),
    to_signed(-1, 8),
    to_signed(-1, 8),
    to_signed(0, 8),
    to_signed(-1, 8),
    to_signed(-1, 8),
    to_signed(-3, 8),
    to_signed(-3, 8),
    to_signed(-3, 8),
    to_signed(-3, 8),
    to_signed(-4, 8),
    to_signed(-4, 8),
    to_signed(-4, 8),
    to_signed(-4, 8),
    to_signed(-3, 8),
    to_signed(-4, 8),
    to_signed(-4, 8),
    to_signed(-5, 8),
    to_signed(-4, 8),
    to_signed(-3, 8),
    to_signed(-3, 8),
    to_signed(-3, 8),
    to_signed(-3, 8),
    to_signed(-3, 8),
    to_signed(-2, 8),
    to_signed(-1, 8),
    to_signed(-1, 8),
    to_signed(-1, 8),
    to_signed(-2, 8),
    to_signed(-2, 8),
    to_signed(-3, 8),
    to_signed(-3, 8),
    to_signed(-3, 8),
    to_signed(-3, 8),
    to_signed(-3, 8),
    to_signed(-3, 8),
    to_signed(-3, 8),
    to_signed(-4, 8),
    to_signed(-4, 8),
    to_signed(-4, 8),
    to_signed(-4, 8),
    to_signed(-4, 8),
    to_signed(-4, 8),
    to_signed(-3, 8),
    to_signed(-4, 8),
    to_signed(-4, 8),
    to_signed(-3, 8),
    to_signed(-2, 8),
    to_signed(-2, 8),
    to_signed(-3, 8),
    to_signed(-4, 8),
    to_signed(-5, 8),
    to_signed(-5, 8),
    to_signed(-5, 8),
    to_signed(-5, 8),
    to_signed(-5, 8),
    to_signed(-6, 8),
    to_signed(-6, 8),
    to_signed(-5, 8),
    to_signed(-5, 8),
    to_signed(-5, 8),
    to_signed(-5, 8),
    to_signed(-5, 8),
    to_signed(-5, 8),
    to_signed(-5, 8),
    to_signed(-4, 8),
    to_signed(-4, 8),
    to_signed(-4, 8),
    to_signed(-4, 8),
    to_signed(-3, 8),
    to_signed(-2, 8),
    to_signed(-3, 8),
    to_signed(-4, 8),
    to_signed(-5, 8),
    to_signed(-5, 8),
    to_signed(-5, 8),
    to_signed(-5, 8),
    to_signed(-5, 8),
    to_signed(-6, 8),
    to_signed(-6, 8),
    to_signed(-6, 8),
    to_signed(-6, 8),
    to_signed(-6, 8),
    to_signed(-6, 8),
    to_signed(-5, 8),
    to_signed(-5, 8),
    to_signed(-5, 8),
    to_signed(-5, 8),
    to_signed(-5, 8),
    to_signed(-5, 8),
    to_signed(-4, 8),
    to_signed(-3, 8),
    to_signed(-2, 8),
    to_signed(-3, 8),
    to_signed(-4, 8),
    to_signed(-5, 8),
    to_signed(-5, 8),
    to_signed(-5, 8),
    to_signed(-4, 8),
    to_signed(-4, 8),
    to_signed(-4, 8),
    to_signed(-4, 8),
    to_signed(-4, 8),
    to_signed(-4, 8),
    to_signed(-3, 8),
    to_signed(-3, 8),
    to_signed(-2, 8),
    to_signed(-1, 8),
    to_signed(-1, 8),
    to_signed(-1, 8),
    to_signed(-1, 8),
    to_signed(-1, 8),
    to_signed(0, 8),
    to_signed(1, 8),
    to_signed(2, 8),
    to_signed(1, 8),
    to_signed(0, 8),
    to_signed(-1, 8),
    to_signed(-2, 8),
    to_signed(-2, 8),
    to_signed(-2, 8),
    to_signed(-1, 8),
    to_signed(-2, 8),
    to_signed(-2, 8),
    to_signed(-2, 8),
    to_signed(-2, 8),
    to_signed(-2, 8),
    to_signed(-1, 8),
    to_signed(-1, 8),
    to_signed(-1, 8),
    to_signed(-2, 8),
    to_signed(-2, 8),
    to_signed(-2, 8),
    to_signed(-2, 8),
    to_signed(-1, 8),
    to_signed(0, 8),
    to_signed(1, 8),
    to_signed(1, 8),
    to_signed(0, 8),
    to_signed(-1, 8),
    to_signed(-2, 8),
    to_signed(-2, 8),
    to_signed(-2, 8),
    to_signed(-2, 8),
    to_signed(-3, 8),
    to_signed(-3, 8),
    to_signed(-3, 8),
    to_signed(-3, 8),
    to_signed(-3, 8),
    to_signed(-3, 8),
    to_signed(-2, 8),
    to_signed(-2, 8),
    to_signed(-3, 8),
    to_signed(-3, 8),
    to_signed(-3, 8),
    to_signed(-2, 8),
    to_signed(-1, 8),
    to_signed(0, 8),
    to_signed(2, 8),
    to_signed(2, 8),
    to_signed(0, 8),
    to_signed(-1, 8),
    to_signed(-2, 8),
    to_signed(-2, 8),
    to_signed(-2, 8),
    to_signed(-2, 8),
    to_signed(-2, 8),
    to_signed(-2, 8),
    to_signed(-2, 8),
    to_signed(-2, 8),
    to_signed(-1, 8),
    to_signed(0, 8),
    to_signed(0, 8),
    to_signed(0, 8),
    to_signed(-1, 8),
    to_signed(-1, 8),
    to_signed(-1, 8),
    to_signed(0, 8),
    to_signed(1, 8),
    to_signed(3, 8),
    to_signed(4, 8),
    to_signed(4, 8),
    to_signed(3, 8),
    to_signed(2, 8),
    to_signed(1, 8),
    to_signed(1, 8),
    to_signed(1, 8),
    to_signed(1, 8),
    to_signed(2, 8),
    to_signed(1, 8),
    to_signed(2, 8),
    to_signed(2, 8),
    to_signed(3, 8),
    to_signed(4, 8),
    to_signed(4, 8),
    to_signed(3, 8),
    to_signed(2, 8),
    to_signed(2, 8),
    to_signed(2, 8),
    to_signed(2, 8),
    to_signed(3, 8),
    to_signed(4, 8),
    to_signed(6, 8),
    to_signed(6, 8),
    to_signed(5, 8),
    to_signed(4, 8),
    to_signed(3, 8),
    to_signed(2, 8),
    to_signed(2, 8),
    to_signed(2, 8),
    to_signed(1, 8),
    to_signed(1, 8),
    to_signed(1, 8),
    to_signed(1, 8),
    to_signed(1, 8),
    to_signed(2, 8),
    to_signed(1, 8),
    to_signed(1, 8),
    to_signed(0, 8),
    to_signed(0, 8),
    to_signed(-1, 8),
    to_signed(-1, 8),
    to_signed(0, 8),
    to_signed(2, 8),
    to_signed(4, 8),
    to_signed(4, 8),
    to_signed(3, 8),
    to_signed(2, 8),
    to_signed(0, 8),
    to_signed(0, 8),
    to_signed(0, 8),
    to_signed(0, 8),
    to_signed(0, 8),
    to_signed(0, 8),
    to_signed(-1, 8),
    to_signed(-1, 8),
    to_signed(0, 8),
    to_signed(1, 8),
    to_signed(2, 8),
    to_signed(1, 8),
    to_signed(0, 8),
    to_signed(0, 8),
    to_signed(0, 8),
    to_signed(0, 8),
    to_signed(1, 8),
    to_signed(4, 8),
    to_signed(5, 8),
    to_signed(6, 8),
    to_signed(5, 8),
    to_signed(4, 8),
    to_signed(3, 8),
    to_signed(3, 8),
    to_signed(3, 8),
    to_signed(3, 8),
    to_signed(3, 8),
    to_signed(2, 8),
    to_signed(2, 8),
    to_signed(2, 8),
    to_signed(2, 8),
    to_signed(3, 8),
    to_signed(3, 8),
    to_signed(2, 8),
    to_signed(0, 8),
    to_signed(0, 8),
    to_signed(-1, 8),
    to_signed(-1, 8),
    to_signed(0, 8),
    to_signed(2, 8),
    to_signed(3, 8),
    to_signed(3, 8),
    to_signed(3, 8),
    to_signed(1, 8),
    to_signed(0, 8),
    to_signed(-1, 8),
    to_signed(-1, 8),
    to_signed(-2, 8),
    to_signed(-2, 8),
    to_signed(-2, 8),
    to_signed(-2, 8),
    to_signed(-1, 8),
    to_signed(-1, 8),
    to_signed(0, 8),
    to_signed(0, 8),
    to_signed(-1, 8),
    to_signed(-2, 8),
    to_signed(-2, 8),
    to_signed(-2, 8),
    to_signed(-2, 8),
    to_signed(-1, 8),
    to_signed(0, 8),
    to_signed(3, 8),
    to_signed(4, 8),
    to_signed(3, 8),
    to_signed(2, 8),
    to_signed(1, 8),
    to_signed(1, 8),
    to_signed(0, 8),
    to_signed(1, 8),
    to_signed(1, 8),
    to_signed(1, 8),
    to_signed(1, 8),
    to_signed(2, 8),
    to_signed(3, 8),
    to_signed(4, 8),
    to_signed(5, 8),
    to_signed(4, 8),
    to_signed(3, 8),
    to_signed(2, 8),
    to_signed(2, 8),
    to_signed(2, 8),
    to_signed(2, 8),
    to_signed(4, 8),
    to_signed(5, 8),
    to_signed(6, 8),
    to_signed(5, 8),
    to_signed(4, 8),
    to_signed(2, 8),
    to_signed(1, 8),
    to_signed(1, 8),
    to_signed(0, 8),
    to_signed(0, 8),
    to_signed(0, 8),
    to_signed(-1, 8),
    to_signed(-1, 8),
    to_signed(0, 8),
    to_signed(1, 8),
    to_signed(1, 8),
    to_signed(0, 8),
    to_signed(-2, 8),
    to_signed(-3, 8),
    to_signed(-3, 8),
    to_signed(-3, 8),
    to_signed(-3, 8),
    to_signed(-1, 8),
    to_signed(0, 8),
    to_signed(1, 8),
    to_signed(1, 8),
    to_signed(0, 8),
    to_signed(-1, 8),
    to_signed(-2, 8),
    to_signed(-2, 8),
    to_signed(-2, 8),
    to_signed(-2, 8),
    to_signed(-2, 8),
    to_signed(-2, 8),
    to_signed(-1, 8),
    to_signed(1, 8),
    to_signed(2, 8),
    to_signed(3, 8),
    to_signed(3, 8),
    to_signed(2, 8),
    to_signed(1, 8),
    to_signed(1, 8),
    to_signed(2, 8),
    to_signed(3, 8),
    to_signed(5, 8),
    to_signed(7, 8),
    to_signed(8, 8),
    to_signed(8, 8),
    to_signed(7, 8),
    to_signed(6, 8),
    to_signed(5, 8),
    to_signed(5, 8),
    to_signed(5, 8),
    to_signed(4, 8),
    to_signed(4, 8),
    to_signed(3, 8),
    to_signed(4, 8),
    to_signed(5, 8),
    to_signed(5, 8),
    to_signed(5, 8),
    to_signed(3, 8),

    to_signed(0, 8)
  );
end package;

